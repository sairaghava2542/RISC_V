 stall_ctrl ( rst, stallreq_if, stallreq_id, stallreq_ex, stallreq_mem, 
        stall );
  output [5:0] stall;
  input rst, stallreq_if, stallreq_id, stallreq_ex, stallreq_mem;
  wire   n3;
  assign stall[3] = stall[4];
  assign stall[0] = stall[1];

  AND2X1_LVT U4 ( .A1(stallreq_mem), .A2(n3), .Y(stall[4]) );
  OA21X1_LVT U5 ( .A1(stallreq_mem), .A2(stallreq_id), .A3(n3), .Y(stall[2])
         );
  AO21X1_LVT U6 ( .A1(stallreq_if), .A2(n3), .A3(stall[2]), .Y(stall[1]) );
  INVX1_LVT U3 ( .A(rst), .Y(n3) );
endmodule


module program_counter ( clk, rst, stall, br, br_addr, pc_o, right_one_o );
  input [5:0] stall;
  input [31:0] br_addr;
  output [31:0] pc_o;
  input clk, rst, br;
  output right_one_o;
  wire   right_one, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n2, n4,
         n6, n8, n9, n11, n46, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n175, n176, n177, n178, n179,
         n181, n182, n183, n184, n185, n186, n188, n189, n191, n192, n193,
         n195, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246;
  wire   [31:0] pc;

  DFFX1_LVT \pc_o_reg[31]  ( .D(n43), .CLK(clk), .Q(pc_o[31]) );
  DFFX1_LVT \pc_o_reg[30]  ( .D(n42), .CLK(clk), .Q(pc_o[30]) );
  DFFX1_LVT \pc_o_reg[29]  ( .D(n41), .CLK(clk), .Q(pc_o[29]) );
  DFFX1_LVT \pc_o_reg[28]  ( .D(n40), .CLK(clk), .Q(pc_o[28]) );
  DFFX1_LVT \pc_o_reg[27]  ( .D(n39), .CLK(clk), .Q(pc_o[27]) );
  DFFX1_LVT \pc_o_reg[26]  ( .D(n38), .CLK(clk), .Q(pc_o[26]) );
  DFFX1_LVT \pc_o_reg[25]  ( .D(n37), .CLK(clk), .Q(pc_o[25]) );
  DFFX1_LVT \pc_o_reg[24]  ( .D(n36), .CLK(clk), .Q(pc_o[24]) );
  DFFX1_LVT \pc_o_reg[23]  ( .D(n35), .CLK(clk), .Q(pc_o[23]) );
  DFFX1_LVT \pc_o_reg[22]  ( .D(n34), .CLK(clk), .Q(pc_o[22]) );
  DFFX1_LVT \pc_o_reg[21]  ( .D(n33), .CLK(clk), .Q(pc_o[21]) );
  DFFX1_LVT \pc_o_reg[20]  ( .D(n32), .CLK(clk), .Q(pc_o[20]) );
  DFFX1_LVT \pc_o_reg[19]  ( .D(n31), .CLK(clk), .Q(pc_o[19]) );
  DFFX1_LVT \pc_o_reg[18]  ( .D(n30), .CLK(clk), .Q(pc_o[18]) );
  DFFX1_LVT \pc_o_reg[17]  ( .D(n29), .CLK(clk), .Q(pc_o[17]) );
  DFFX1_LVT \pc_o_reg[16]  ( .D(n28), .CLK(clk), .Q(pc_o[16]) );
  DFFX1_LVT \pc_o_reg[15]  ( .D(n27), .CLK(clk), .Q(pc_o[15]) );
  DFFX1_LVT \pc_o_reg[14]  ( .D(n26), .CLK(clk), .Q(pc_o[14]) );
  DFFX1_LVT \pc_o_reg[13]  ( .D(n25), .CLK(clk), .Q(pc_o[13]) );
  DFFX1_LVT \pc_o_reg[12]  ( .D(n24), .CLK(clk), .Q(pc_o[12]) );
  DFFX1_LVT \pc_o_reg[11]  ( .D(n23), .CLK(clk), .Q(pc_o[11]) );
  DFFX1_LVT \pc_o_reg[10]  ( .D(n22), .CLK(clk), .Q(pc_o[10]) );
  DFFX1_LVT \pc_o_reg[9]  ( .D(n21), .CLK(clk), .Q(pc_o[9]) );
  DFFX1_LVT \pc_o_reg[8]  ( .D(n20), .CLK(clk), .Q(pc_o[8]) );
  DFFX1_LVT \pc_o_reg[7]  ( .D(n19), .CLK(clk), .Q(pc_o[7]) );
  DFFX1_LVT \pc_o_reg[6]  ( .D(n18), .CLK(clk), .Q(pc_o[6]) );
  DFFX1_LVT \pc_o_reg[5]  ( .D(n17), .CLK(clk), .Q(pc_o[5]) );
  DFFX1_LVT \pc_o_reg[4]  ( .D(n16), .CLK(clk), .Q(pc_o[4]) );
  DFFX1_LVT \pc_o_reg[3]  ( .D(n15), .CLK(clk), .Q(pc_o[3]) );
  DFFX1_LVT \pc_o_reg[2]  ( .D(n14), .CLK(clk), .Q(pc_o[2]) );
  DFFX1_LVT \pc_o_reg[1]  ( .D(n13), .CLK(clk), .Q(pc_o[1]) );
  DFFX1_LVT \pc_o_reg[0]  ( .D(n12), .CLK(clk), .Q(pc_o[0]) );
  DFFX1_LVT right_one_o_reg ( .D(n44), .CLK(clk), .Q(right_one_o) );
  DFFX1_LVT right_one_reg ( .D(n45), .CLK(clk), .Q(right_one) );
  DFFX1_LVT \pc_reg[1]  ( .D(n77), .CLK(clk), .Q(pc[1]) );
  DFFX1_LVT \pc_reg[0]  ( .D(n78), .CLK(clk), .Q(pc[0]) );
  DFFX1_LVT \pc_reg[31]  ( .D(n47), .CLK(clk), .Q(pc[31]), .QN(n233) );
  DFFX1_LVT \pc_reg[30]  ( .D(n48), .CLK(clk), .Q(pc[30]), .QN(n232) );
  DFFX1_LVT \pc_reg[26]  ( .D(n52), .CLK(clk), .Q(pc[26]), .QN(n228) );
  DFFX1_LVT \pc_reg[24]  ( .D(n54), .CLK(clk), .Q(pc[24]), .QN(n226) );
  DFFX1_LVT \pc_reg[22]  ( .D(n56), .CLK(clk), .Q(pc[22]), .QN(n224) );
  DFFX1_LVT \pc_reg[18]  ( .D(n60), .CLK(clk), .Q(pc[18]), .QN(n220) );
  DFFX1_LVT \pc_reg[16]  ( .D(n62), .CLK(clk), .Q(pc[16]), .QN(n218) );
  OA221X1_LVT U5 ( .A1(br), .A2(pc[0]), .A3(n235), .A4(br_addr[0]), .A5(n234), 
        .Y(n78) );
  OA221X1_LVT U6 ( .A1(br), .A2(pc[1]), .A3(n235), .A4(br_addr[1]), .A5(n234), 
        .Y(n77) );
  NAND2X0_LVT U10 ( .A1(br), .A2(n234), .Y(n8) );
  AOI22X1_LVT U13 ( .A1(br), .A2(br_addr[2]), .A3(pc[2]), .A4(n238), .Y(n6) );
  NAND2X0_LVT U18 ( .A1(n237), .A2(n8), .Y(n81) );
  NAND2X0_LVT U21 ( .A1(n240), .A2(n204), .Y(n4) );
  NAND3X0_LVT U22 ( .A1(n6), .A2(n234), .A3(n4), .Y(n76) );
  AO21X1_LVT U24 ( .A1(n204), .A2(n240), .A3(n238), .Y(n11) );
  AND2X1_LVT U25 ( .A1(n240), .A2(n206), .Y(n9) );
  AO222X1_LVT U28 ( .A1(n11), .A2(pc[3]), .A3(pc[2]), .A4(n9), .A5(n236), .A6(
        br_addr[3]), .Y(n75) );
  NAND4X0_LVT U29 ( .A1(n240), .A2(pc[2]), .A3(pc[3]), .A4(n205), .Y(n80) );
  NAND2X0_LVT U31 ( .A1(br_addr[4]), .A2(n236), .Y(n79) );
  OAI221X1_LVT U32 ( .A1(n11), .A2(n206), .A3(n11), .A4(n240), .A5(pc[4]), .Y(
        n46) );
  NAND3X0_LVT U33 ( .A1(n80), .A2(n79), .A3(n46), .Y(n74) );
  AND3X1_LVT U34 ( .A1(pc[4]), .A2(pc[2]), .A3(pc[3]), .Y(n89) );
  OA21X1_LVT U36 ( .A1(n89), .A2(n239), .A3(n179), .Y(n85) );
  NAND2X0_LVT U37 ( .A1(n240), .A2(n89), .Y(n82) );
  AO22X1_LVT U38 ( .A1(pc[5]), .A2(n85), .A3(n207), .A4(n82), .Y(n84) );
  NAND2X0_LVT U39 ( .A1(n236), .A2(br_addr[5]), .Y(n83) );
  NAND2X0_LVT U40 ( .A1(n84), .A2(n83), .Y(n73) );
  NAND4X0_LVT U41 ( .A1(pc[5]), .A2(n240), .A3(n89), .A4(n208), .Y(n88) );
  NAND2X0_LVT U42 ( .A1(br_addr[6]), .A2(n236), .Y(n87) );
  AO221X1_LVT U43 ( .A1(n85), .A2(pc[5]), .A3(n85), .A4(n239), .A5(n208), .Y(
        n86) );
  NAND3X0_LVT U44 ( .A1(n88), .A2(n87), .A3(n86), .Y(n72) );
  AND3X1_LVT U45 ( .A1(pc[5]), .A2(pc[6]), .A3(n89), .Y(n97) );
  OA21X1_LVT U46 ( .A1(n97), .A2(n239), .A3(n179), .Y(n93) );
  NAND2X0_LVT U47 ( .A1(n240), .A2(n97), .Y(n90) );
  AO22X1_LVT U48 ( .A1(n244), .A2(n93), .A3(n209), .A4(n90), .Y(n92) );
  NAND2X0_LVT U49 ( .A1(n236), .A2(br_addr[7]), .Y(n91) );
  NAND2X0_LVT U50 ( .A1(n92), .A2(n91), .Y(n71) );
  NAND4X0_LVT U51 ( .A1(n244), .A2(n240), .A3(n97), .A4(n210), .Y(n96) );
  NAND2X0_LVT U52 ( .A1(br_addr[8]), .A2(n236), .Y(n95) );
  AO221X1_LVT U53 ( .A1(n93), .A2(pc[7]), .A3(n93), .A4(n239), .A5(n210), .Y(
        n94) );
  NAND3X0_LVT U54 ( .A1(n96), .A2(n95), .A3(n94), .Y(n70) );
  AND3X1_LVT U55 ( .A1(pc[7]), .A2(pc[8]), .A3(n97), .Y(n105) );
  OA21X1_LVT U56 ( .A1(n105), .A2(n239), .A3(n179), .Y(n101) );
  NAND2X0_LVT U57 ( .A1(n240), .A2(n105), .Y(n98) );
  AO22X1_LVT U58 ( .A1(n245), .A2(n101), .A3(n211), .A4(n98), .Y(n100) );
  NAND2X0_LVT U59 ( .A1(n236), .A2(br_addr[9]), .Y(n99) );
  NAND2X0_LVT U60 ( .A1(n100), .A2(n99), .Y(n69) );
  NAND4X0_LVT U61 ( .A1(n245), .A2(n240), .A3(n105), .A4(n212), .Y(n104) );
  NAND2X0_LVT U62 ( .A1(br_addr[10]), .A2(n236), .Y(n103) );
  AO221X1_LVT U63 ( .A1(n101), .A2(pc[9]), .A3(n101), .A4(n239), .A5(n212), 
        .Y(n102) );
  NAND3X0_LVT U64 ( .A1(n104), .A2(n103), .A3(n102), .Y(n68) );
  AND3X1_LVT U65 ( .A1(pc[9]), .A2(pc[10]), .A3(n105), .Y(n113) );
  OA21X1_LVT U66 ( .A1(n113), .A2(n239), .A3(n179), .Y(n109) );
  NAND2X0_LVT U67 ( .A1(n240), .A2(n113), .Y(n106) );
  AO22X1_LVT U68 ( .A1(n243), .A2(n109), .A3(n213), .A4(n106), .Y(n108) );
  NAND2X0_LVT U69 ( .A1(n236), .A2(br_addr[11]), .Y(n107) );
  NAND2X0_LVT U70 ( .A1(n108), .A2(n107), .Y(n67) );
  NAND4X0_LVT U71 ( .A1(n243), .A2(n240), .A3(n113), .A4(n214), .Y(n112) );
  NAND2X0_LVT U72 ( .A1(br_addr[12]), .A2(n236), .Y(n111) );
  AO221X1_LVT U73 ( .A1(n109), .A2(n243), .A3(n109), .A4(n239), .A5(n214), .Y(
        n110) );
  NAND3X0_LVT U74 ( .A1(n112), .A2(n111), .A3(n110), .Y(n66) );
  AND3X1_LVT U75 ( .A1(pc[11]), .A2(pc[12]), .A3(n113), .Y(n121) );
  OA21X1_LVT U76 ( .A1(n121), .A2(n241), .A3(n179), .Y(n117) );
  NAND2X0_LVT U77 ( .A1(n242), .A2(n121), .Y(n114) );
  AO22X1_LVT U78 ( .A1(pc[13]), .A2(n117), .A3(n215), .A4(n114), .Y(n116) );
  NAND2X0_LVT U79 ( .A1(n236), .A2(br_addr[13]), .Y(n115) );
  NAND2X0_LVT U80 ( .A1(n116), .A2(n115), .Y(n65) );
  NAND4X0_LVT U81 ( .A1(pc[13]), .A2(n242), .A3(n121), .A4(n216), .Y(n120) );
  NAND2X0_LVT U82 ( .A1(br_addr[14]), .A2(n236), .Y(n119) );
  AO221X1_LVT U83 ( .A1(n117), .A2(pc[13]), .A3(n117), .A4(n241), .A5(n216), 
        .Y(n118) );
  NAND3X0_LVT U84 ( .A1(n120), .A2(n119), .A3(n118), .Y(n64) );
  AND3X1_LVT U85 ( .A1(pc[13]), .A2(pc[14]), .A3(n121), .Y(n129) );
  OA21X1_LVT U86 ( .A1(n129), .A2(n241), .A3(n179), .Y(n125) );
  NAND2X0_LVT U87 ( .A1(n242), .A2(n129), .Y(n122) );
  AO22X1_LVT U88 ( .A1(pc[15]), .A2(n125), .A3(n217), .A4(n122), .Y(n124) );
  NAND2X0_LVT U89 ( .A1(n236), .A2(br_addr[15]), .Y(n123) );
  NAND2X0_LVT U90 ( .A1(n124), .A2(n123), .Y(n63) );
  NAND4X0_LVT U91 ( .A1(pc[15]), .A2(n242), .A3(n129), .A4(n218), .Y(n128) );
  NAND2X0_LVT U92 ( .A1(br_addr[16]), .A2(n236), .Y(n127) );
  AO221X1_LVT U93 ( .A1(n125), .A2(pc[15]), .A3(n125), .A4(n241), .A5(n218), 
        .Y(n126) );
  NAND3X0_LVT U94 ( .A1(n128), .A2(n127), .A3(n126), .Y(n62) );
  AND3X1_LVT U95 ( .A1(pc[15]), .A2(pc[16]), .A3(n129), .Y(n137) );
  OA21X1_LVT U96 ( .A1(n137), .A2(n241), .A3(n179), .Y(n133) );
  NAND2X0_LVT U97 ( .A1(n242), .A2(n137), .Y(n130) );
  AO22X1_LVT U98 ( .A1(pc[17]), .A2(n133), .A3(n219), .A4(n130), .Y(n132) );
  NAND2X0_LVT U99 ( .A1(n236), .A2(br_addr[17]), .Y(n131) );
  NAND2X0_LVT U100 ( .A1(n132), .A2(n131), .Y(n61) );
  NAND4X0_LVT U101 ( .A1(pc[17]), .A2(n242), .A3(n137), .A4(n220), .Y(n136) );
  NAND2X0_LVT U102 ( .A1(br_addr[18]), .A2(n236), .Y(n135) );
  AO221X1_LVT U103 ( .A1(n133), .A2(pc[17]), .A3(n133), .A4(n241), .A5(n220), 
        .Y(n134) );
  NAND3X0_LVT U104 ( .A1(n136), .A2(n135), .A3(n134), .Y(n60) );
  AND3X1_LVT U105 ( .A1(pc[17]), .A2(pc[18]), .A3(n137), .Y(n145) );
  OA21X1_LVT U106 ( .A1(n145), .A2(n241), .A3(n179), .Y(n141) );
  NAND2X0_LVT U107 ( .A1(n242), .A2(n145), .Y(n138) );
  AO22X1_LVT U108 ( .A1(pc[19]), .A2(n141), .A3(n221), .A4(n138), .Y(n140) );
  NAND2X0_LVT U109 ( .A1(n236), .A2(br_addr[19]), .Y(n139) );
  NAND2X0_LVT U110 ( .A1(n140), .A2(n139), .Y(n59) );
  NAND4X0_LVT U111 ( .A1(pc[19]), .A2(n242), .A3(n145), .A4(n222), .Y(n144) );
  NAND2X0_LVT U112 ( .A1(br_addr[20]), .A2(n236), .Y(n143) );
  AO221X1_LVT U113 ( .A1(n141), .A2(pc[19]), .A3(n141), .A4(n241), .A5(n222), 
        .Y(n142) );
  NAND3X0_LVT U114 ( .A1(n144), .A2(n143), .A3(n142), .Y(n58) );
  AND3X1_LVT U115 ( .A1(pc[19]), .A2(pc[20]), .A3(n145), .Y(n153) );
  OA21X1_LVT U116 ( .A1(n153), .A2(n239), .A3(n179), .Y(n149) );
  NAND2X0_LVT U117 ( .A1(n240), .A2(n153), .Y(n146) );
  AO22X1_LVT U118 ( .A1(pc[21]), .A2(n149), .A3(n223), .A4(n146), .Y(n148) );
  NAND2X0_LVT U119 ( .A1(n236), .A2(br_addr[21]), .Y(n147) );
  NAND2X0_LVT U120 ( .A1(n148), .A2(n147), .Y(n57) );
  NAND4X0_LVT U121 ( .A1(pc[21]), .A2(n240), .A3(n153), .A4(n224), .Y(n152) );
  NAND2X0_LVT U122 ( .A1(br_addr[22]), .A2(n236), .Y(n151) );
  AO221X1_LVT U123 ( .A1(n149), .A2(pc[21]), .A3(n149), .A4(n239), .A5(n224), 
        .Y(n150) );
  NAND3X0_LVT U124 ( .A1(n152), .A2(n151), .A3(n150), .Y(n56) );
  AND3X1_LVT U125 ( .A1(pc[21]), .A2(pc[22]), .A3(n153), .Y(n161) );
  OA21X1_LVT U126 ( .A1(n161), .A2(n239), .A3(n179), .Y(n157) );
  NAND2X0_LVT U127 ( .A1(n240), .A2(n161), .Y(n154) );
  AO22X1_LVT U128 ( .A1(pc[23]), .A2(n157), .A3(n225), .A4(n154), .Y(n156) );
  NAND2X0_LVT U129 ( .A1(n236), .A2(br_addr[23]), .Y(n155) );
  NAND2X0_LVT U130 ( .A1(n156), .A2(n155), .Y(n55) );
  NAND4X0_LVT U131 ( .A1(pc[23]), .A2(n240), .A3(n161), .A4(n226), .Y(n160) );
  NAND2X0_LVT U132 ( .A1(br_addr[24]), .A2(n236), .Y(n159) );
  AO221X1_LVT U133 ( .A1(n157), .A2(pc[23]), .A3(n157), .A4(n239), .A5(n226), 
        .Y(n158) );
  NAND3X0_LVT U134 ( .A1(n160), .A2(n159), .A3(n158), .Y(n54) );
  AND3X1_LVT U135 ( .A1(pc[23]), .A2(pc[24]), .A3(n161), .Y(n169) );
  OA21X1_LVT U136 ( .A1(n169), .A2(n239), .A3(n179), .Y(n165) );
  NAND2X0_LVT U137 ( .A1(n240), .A2(n169), .Y(n162) );
  AO22X1_LVT U138 ( .A1(pc[25]), .A2(n165), .A3(n227), .A4(n162), .Y(n164) );
  NAND2X0_LVT U139 ( .A1(n236), .A2(br_addr[25]), .Y(n163) );
  NAND2X0_LVT U140 ( .A1(n164), .A2(n163), .Y(n53) );
  NAND4X0_LVT U141 ( .A1(pc[25]), .A2(n240), .A3(n169), .A4(n228), .Y(n168) );
  NAND2X0_LVT U142 ( .A1(br_addr[26]), .A2(n236), .Y(n167) );
  AO221X1_LVT U143 ( .A1(n165), .A2(pc[25]), .A3(n165), .A4(n239), .A5(n228), 
        .Y(n166) );
  NAND3X0_LVT U144 ( .A1(n168), .A2(n167), .A3(n166), .Y(n52) );
  AND3X1_LVT U145 ( .A1(pc[25]), .A2(pc[26]), .A3(n169), .Y(n182) );
  OA21X1_LVT U146 ( .A1(n182), .A2(n241), .A3(n179), .Y(n175) );
  NAND2X0_LVT U147 ( .A1(n242), .A2(n182), .Y(n170) );
  AO22X1_LVT U148 ( .A1(pc[27]), .A2(n175), .A3(n229), .A4(n170), .Y(n172) );
  NAND2X0_LVT U149 ( .A1(n236), .A2(br_addr[27]), .Y(n171) );
  NAND2X0_LVT U150 ( .A1(n172), .A2(n171), .Y(n51) );
  NAND4X0_LVT U151 ( .A1(pc[27]), .A2(n242), .A3(n182), .A4(n230), .Y(n178) );
  NAND2X0_LVT U152 ( .A1(br_addr[28]), .A2(n236), .Y(n177) );
  AO221X1_LVT U153 ( .A1(n175), .A2(pc[27]), .A3(n175), .A4(n241), .A5(n230), 
        .Y(n176) );
  NAND3X0_LVT U154 ( .A1(n178), .A2(n177), .A3(n176), .Y(n50) );
  AND3X1_LVT U155 ( .A1(pc[27]), .A2(pc[28]), .A3(n182), .Y(n181) );
  OAI21X1_LVT U156 ( .A1(n181), .A2(n241), .A3(n179), .Y(n184) );
  AND4X1_LVT U157 ( .A1(n242), .A2(pc[27]), .A3(pc[28]), .A4(n182), .Y(n185)
         );
  AO22X1_LVT U158 ( .A1(n236), .A2(br_addr[29]), .A3(n185), .A4(n231), .Y(n183) );
  AO21X1_LVT U159 ( .A1(pc[29]), .A2(n184), .A3(n183), .Y(n49) );
  AO21X1_LVT U160 ( .A1(n231), .A2(n242), .A3(n184), .Y(n188) );
  AND2X1_LVT U161 ( .A1(pc[29]), .A2(n185), .Y(n189) );
  AO22X1_LVT U162 ( .A1(br_addr[30]), .A2(n236), .A3(n189), .A4(n232), .Y(n186) );
  AO21X1_LVT U163 ( .A1(pc[30]), .A2(n188), .A3(n186), .Y(n48) );
  OAI221X1_LVT U164 ( .A1(n188), .A2(n232), .A3(n188), .A4(n242), .A5(pc[31]), 
        .Y(n193) );
  NAND3X0_LVT U165 ( .A1(pc[30]), .A2(n189), .A3(n233), .Y(n192) );
  NAND2X0_LVT U166 ( .A1(br_addr[31]), .A2(n236), .Y(n191) );
  NAND3X0_LVT U167 ( .A1(n193), .A2(n192), .A3(n191), .Y(n47) );
  AO21X1_LVT U168 ( .A1(n2), .A2(right_one), .A3(n236), .Y(n45) );
  AO22X1_LVT U169 ( .A1(n237), .A2(right_one), .A3(n195), .A4(right_one_o), 
        .Y(n44) );
  AO22X1_LVT U171 ( .A1(pc[31]), .A2(n237), .A3(n246), .A4(pc_o[31]), .Y(n43)
         );
  AO22X1_LVT U172 ( .A1(pc[30]), .A2(n237), .A3(n246), .A4(pc_o[30]), .Y(n42)
         );
  AO22X1_LVT U174 ( .A1(n237), .A2(pc[29]), .A3(n246), .A4(pc_o[29]), .Y(n41)
         );
  AO22X1_LVT U176 ( .A1(n237), .A2(pc[28]), .A3(n246), .A4(pc_o[28]), .Y(n40)
         );
  AO22X1_LVT U177 ( .A1(n237), .A2(pc[27]), .A3(n2), .A4(pc_o[27]), .Y(n39) );
  AO22X1_LVT U178 ( .A1(n237), .A2(pc[26]), .A3(n246), .A4(pc_o[26]), .Y(n38)
         );
  AO22X1_LVT U179 ( .A1(n237), .A2(pc[25]), .A3(n246), .A4(pc_o[25]), .Y(n37)
         );
  AO22X1_LVT U180 ( .A1(n237), .A2(pc[24]), .A3(n2), .A4(pc_o[24]), .Y(n36) );
  AO22X1_LVT U181 ( .A1(n237), .A2(pc[23]), .A3(n246), .A4(pc_o[23]), .Y(n35)
         );
  AO22X1_LVT U182 ( .A1(n237), .A2(pc[22]), .A3(n246), .A4(pc_o[22]), .Y(n34)
         );
  AO22X1_LVT U183 ( .A1(n237), .A2(pc[21]), .A3(n246), .A4(pc_o[21]), .Y(n33)
         );
  AO22X1_LVT U184 ( .A1(n237), .A2(pc[20]), .A3(n246), .A4(pc_o[20]), .Y(n32)
         );
  AO22X1_LVT U185 ( .A1(n237), .A2(pc[19]), .A3(n246), .A4(pc_o[19]), .Y(n31)
         );
  AO22X1_LVT U186 ( .A1(n237), .A2(pc[18]), .A3(n246), .A4(pc_o[18]), .Y(n30)
         );
  AO22X1_LVT U187 ( .A1(n237), .A2(pc[17]), .A3(n246), .A4(pc_o[17]), .Y(n29)
         );
  AO22X1_LVT U188 ( .A1(n237), .A2(pc[16]), .A3(n246), .A4(pc_o[16]), .Y(n28)
         );
  AO22X1_LVT U189 ( .A1(n237), .A2(pc[15]), .A3(n246), .A4(pc_o[15]), .Y(n27)
         );
  AO22X1_LVT U191 ( .A1(n237), .A2(pc[14]), .A3(n246), .A4(pc_o[14]), .Y(n26)
         );
  AO22X1_LVT U192 ( .A1(n237), .A2(pc[13]), .A3(n246), .A4(pc_o[13]), .Y(n25)
         );
  AO22X1_LVT U193 ( .A1(n237), .A2(pc[12]), .A3(n246), .A4(pc_o[12]), .Y(n24)
         );
  AO22X1_LVT U194 ( .A1(n237), .A2(n243), .A3(n246), .A4(pc_o[11]), .Y(n23) );
  AO22X1_LVT U195 ( .A1(n237), .A2(pc[10]), .A3(n246), .A4(pc_o[10]), .Y(n22)
         );
  AO22X1_LVT U196 ( .A1(n237), .A2(n245), .A3(n246), .A4(pc_o[9]), .Y(n21) );
  AO22X1_LVT U197 ( .A1(n237), .A2(pc[8]), .A3(n2), .A4(pc_o[8]), .Y(n20) );
  AO22X1_LVT U198 ( .A1(n237), .A2(n244), .A3(n246), .A4(pc_o[7]), .Y(n19) );
  AO22X1_LVT U199 ( .A1(n237), .A2(pc[6]), .A3(n246), .A4(pc_o[6]), .Y(n18) );
  AO22X1_LVT U200 ( .A1(n237), .A2(pc[5]), .A3(n246), .A4(pc_o[5]), .Y(n17) );
  AO22X1_LVT U201 ( .A1(n237), .A2(pc[4]), .A3(n2), .A4(pc_o[4]), .Y(n16) );
  AO22X1_LVT U202 ( .A1(n237), .A2(pc[3]), .A3(n246), .A4(pc_o[3]), .Y(n15) );
  AO22X1_LVT U203 ( .A1(n237), .A2(pc[2]), .A3(n246), .A4(pc_o[2]), .Y(n14) );
  AO22X1_LVT U204 ( .A1(n237), .A2(pc[1]), .A3(n246), .A4(pc_o[1]), .Y(n13) );
  AO22X1_LVT U205 ( .A1(n237), .A2(pc[0]), .A3(n246), .A4(pc_o[0]), .Y(n12) );
  NAND2X2_LVT U11 ( .A1(n2), .A2(n8), .Y(n179) );
  INVX1_LVT U3 ( .A(rst), .Y(n234) );
  INVX1_LVT U4 ( .A(br), .Y(n235) );
  INVX4_LVT U8 ( .A(n8), .Y(n236) );
  INVX8_LVT U9 ( .A(n195), .Y(n237) );
  INVX1_LVT U12 ( .A(n179), .Y(n238) );
  NBUFFX4_LVT U15 ( .A(n81), .Y(n239) );
  INVX2_LVT U16 ( .A(n239), .Y(n240) );
  NBUFFX4_LVT U17 ( .A(n81), .Y(n241) );
  INVX2_LVT U19 ( .A(n241), .Y(n242) );
  AND2X4_LVT U7 ( .A1(stall[0]), .A2(n234), .Y(n2) );
  DFFX2_LVT \pc_reg[5]  ( .D(n73), .CLK(clk), .Q(pc[5]), .QN(n207) );
  DFFX2_LVT \pc_reg[13]  ( .D(n65), .CLK(clk), .Q(pc[13]), .QN(n215) );
  DFFX2_LVT \pc_reg[10]  ( .D(n68), .CLK(clk), .Q(pc[10]), .QN(n212) );
  DFFX2_LVT \pc_reg[8]  ( .D(n70), .CLK(clk), .Q(pc[8]), .QN(n210) );
  DFFX2_LVT \pc_reg[2]  ( .D(n76), .CLK(clk), .Q(pc[2]), .QN(n204) );
  DFFX2_LVT \pc_reg[4]  ( .D(n74), .CLK(clk), .Q(pc[4]), .QN(n205) );
  DFFX2_LVT \pc_reg[3]  ( .D(n75), .CLK(clk), .Q(pc[3]), .QN(n206) );
  DFFX2_LVT \pc_reg[6]  ( .D(n72), .CLK(clk), .Q(pc[6]), .QN(n208) );
  DFFX2_LVT \pc_reg[12]  ( .D(n66), .CLK(clk), .Q(pc[12]), .QN(n214) );
  DFFX2_LVT \pc_reg[17]  ( .D(n61), .CLK(clk), .Q(pc[17]), .QN(n219) );
  DFFX2_LVT \pc_reg[15]  ( .D(n63), .CLK(clk), .Q(pc[15]), .QN(n217) );
  DFFX2_LVT \pc_reg[19]  ( .D(n59), .CLK(clk), .Q(pc[19]), .QN(n221) );
  DFFX2_LVT \pc_reg[27]  ( .D(n51), .CLK(clk), .Q(pc[27]), .QN(n229) );
  DFFX2_LVT \pc_reg[25]  ( .D(n53), .CLK(clk), .Q(pc[25]), .QN(n227) );
  DFFX2_LVT \pc_reg[21]  ( .D(n57), .CLK(clk), .Q(pc[21]), .QN(n223) );
  DFFX2_LVT \pc_reg[14]  ( .D(n64), .CLK(clk), .Q(pc[14]), .QN(n216) );
  OR2X2_LVT U14 ( .A1(stall[0]), .A2(rst), .Y(n195) );
  DFFX2_LVT \pc_reg[23]  ( .D(n55), .CLK(clk), .Q(pc[23]), .QN(n225) );
  DFFX2_LVT \pc_reg[28]  ( .D(n50), .CLK(clk), .Q(pc[28]), .QN(n230) );
  DFFX2_LVT \pc_reg[29]  ( .D(n49), .CLK(clk), .Q(pc[29]), .QN(n231) );
  DFFX2_LVT \pc_reg[20]  ( .D(n58), .CLK(clk), .Q(pc[20]), .QN(n222) );
  DFFX1_LVT \pc_reg[7]  ( .D(n71), .CLK(clk), .Q(pc[7]), .QN(n209) );
  DFFX1_LVT \pc_reg[9]  ( .D(n69), .CLK(clk), .Q(pc[9]), .QN(n211) );
  DFFX1_LVT \pc_reg[11]  ( .D(n67), .CLK(clk), .Q(pc[11]), .QN(n213) );
  NBUFFX4_LVT U20 ( .A(pc[7]), .Y(n244) );
  NBUFFX4_LVT U23 ( .A(pc[11]), .Y(n243) );
  NBUFFX4_LVT U26 ( .A(pc[9]), .Y(n245) );
  NBUFFX4_LVT U27 ( .A(n2), .Y(n246) );
endmodule


module inst_fetch ( rst, pc_i, mem_data_i, mem_busy, mem_done, br, right_one, 
        mem_re, mem_addr_o, pc_o, inst_o, stallreq );
  input [31:0] pc_i;
  input [31:0] mem_data_i;
  input [1:0] mem_busy;
  input [1:0] mem_done;
  output [31:0] mem_addr_o;
  output [31:0] pc_o;
  output [31:0] inst_o;
  input rst, br, right_one;
  output mem_re, stallreq;
  wire   mem_taking, waiting_one, N14, N15, N16, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96,
         N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108,
         N109, N110, N111, N112, N113, N114, N115, N116, N118, N119, n1, n2,
         n5, n6, n9, n12, n13, n14, n15, n24, n35, n36, n37, n38, n39, n40,
         n41, n42, n43;

  LATCHX1_LVT waiting_one_reg ( .CLK(N118), .D(N119), .Q(waiting_one) );
  LATCHX1_LVT \pc_o_reg[0]  ( .CLK(n40), .D(N19), .Q(pc_o[0]) );
  LATCHX1_LVT \inst_o_reg[31]  ( .CLK(n39), .D(N82), .Q(inst_o[31]) );
  LATCHX1_LVT \inst_o_reg[30]  ( .CLK(n39), .D(N81), .Q(inst_o[30]) );
  LATCHX1_LVT \inst_o_reg[29]  ( .CLK(n39), .D(N80), .Q(inst_o[29]) );
  LATCHX1_LVT \inst_o_reg[28]  ( .CLK(n39), .D(N79), .Q(inst_o[28]) );
  LATCHX1_LVT \inst_o_reg[27]  ( .CLK(n39), .D(N78), .Q(inst_o[27]) );
  LATCHX1_LVT \inst_o_reg[26]  ( .CLK(n39), .D(N77), .Q(inst_o[26]) );
  LATCHX1_LVT \inst_o_reg[25]  ( .CLK(n39), .D(N76), .Q(inst_o[25]) );
  LATCHX1_LVT \inst_o_reg[24]  ( .CLK(n39), .D(N75), .Q(inst_o[24]) );
  LATCHX1_LVT \inst_o_reg[23]  ( .CLK(n39), .D(N74), .Q(inst_o[23]) );
  LATCHX1_LVT \inst_o_reg[22]  ( .CLK(n39), .D(N73), .Q(inst_o[22]) );
  LATCHX1_LVT \inst_o_reg[21]  ( .CLK(n39), .D(N72), .Q(inst_o[21]) );
  LATCHX1_LVT \inst_o_reg[20]  ( .CLK(n39), .D(N71), .Q(inst_o[20]) );
  LATCHX1_LVT \inst_o_reg[19]  ( .CLK(n39), .D(N70), .Q(inst_o[19]) );
  LATCHX1_LVT \inst_o_reg[18]  ( .CLK(n39), .D(N69), .Q(inst_o[18]) );
  LATCHX1_LVT \inst_o_reg[17]  ( .CLK(n39), .D(N68), .Q(inst_o[17]) );
  LATCHX1_LVT \inst_o_reg[16]  ( .CLK(n39), .D(N67), .Q(inst_o[16]) );
  LATCHX1_LVT \inst_o_reg[15]  ( .CLK(n39), .D(N66), .Q(inst_o[15]) );
  LATCHX1_LVT \inst_o_reg[14]  ( .CLK(n39), .D(N65), .Q(inst_o[14]) );
  LATCHX1_LVT \inst_o_reg[13]  ( .CLK(n39), .D(N64), .Q(inst_o[13]) );
  LATCHX1_LVT \inst_o_reg[12]  ( .CLK(n39), .D(N63), .Q(inst_o[12]) );
  LATCHX1_LVT \inst_o_reg[11]  ( .CLK(n39), .D(N62), .Q(inst_o[11]) );
  LATCHX1_LVT \inst_o_reg[10]  ( .CLK(n39), .D(N61), .Q(inst_o[10]) );
  LATCHX1_LVT \inst_o_reg[9]  ( .CLK(n39), .D(N60), .Q(inst_o[9]) );
  LATCHX1_LVT \inst_o_reg[8]  ( .CLK(n39), .D(N59), .Q(inst_o[8]) );
  LATCHX1_LVT \inst_o_reg[7]  ( .CLK(n39), .D(N58), .Q(inst_o[7]) );
  LATCHX1_LVT \inst_o_reg[6]  ( .CLK(n39), .D(N57), .Q(inst_o[6]) );
  LATCHX1_LVT \inst_o_reg[5]  ( .CLK(n39), .D(N56), .Q(inst_o[5]) );
  LATCHX1_LVT \inst_o_reg[4]  ( .CLK(n39), .D(N55), .Q(inst_o[4]) );
  LATCHX1_LVT \inst_o_reg[3]  ( .CLK(n39), .D(N54), .Q(inst_o[3]) );
  LATCHX1_LVT \inst_o_reg[2]  ( .CLK(n39), .D(N53), .Q(inst_o[2]) );
  LATCHX1_LVT \inst_o_reg[1]  ( .CLK(n39), .D(N52), .Q(inst_o[1]) );
  LATCHX1_LVT \inst_o_reg[0]  ( .CLK(n39), .D(N51), .Q(inst_o[0]) );
  LATCHX1_LVT \pc_o_reg[31]  ( .CLK(n40), .D(N50), .Q(pc_o[31]) );
  LATCHX1_LVT \pc_o_reg[30]  ( .CLK(n40), .D(N49), .Q(pc_o[30]) );
  LATCHX1_LVT \pc_o_reg[29]  ( .CLK(n40), .D(N48), .Q(pc_o[29]) );
  LATCHX1_LVT \pc_o_reg[28]  ( .CLK(n40), .D(N47), .Q(pc_o[28]) );
  LATCHX1_LVT \pc_o_reg[27]  ( .CLK(n40), .D(N46), .Q(pc_o[27]) );
  LATCHX1_LVT \pc_o_reg[26]  ( .CLK(n40), .D(N45), .Q(pc_o[26]) );
  LATCHX1_LVT \pc_o_reg[25]  ( .CLK(n40), .D(N44), .Q(pc_o[25]) );
  LATCHX1_LVT \pc_o_reg[24]  ( .CLK(n40), .D(N43), .Q(pc_o[24]) );
  LATCHX1_LVT \pc_o_reg[23]  ( .CLK(n40), .D(N42), .Q(pc_o[23]) );
  LATCHX1_LVT \pc_o_reg[22]  ( .CLK(n40), .D(N41), .Q(pc_o[22]) );
  LATCHX1_LVT \pc_o_reg[21]  ( .CLK(n40), .D(N40), .Q(pc_o[21]) );
  LATCHX1_LVT \pc_o_reg[20]  ( .CLK(n40), .D(N39), .Q(pc_o[20]) );
  LATCHX1_LVT \pc_o_reg[19]  ( .CLK(n40), .D(N38), .Q(pc_o[19]) );
  LATCHX1_LVT \pc_o_reg[18]  ( .CLK(n40), .D(N37), .Q(pc_o[18]) );
  LATCHX1_LVT \pc_o_reg[17]  ( .CLK(n40), .D(N36), .Q(pc_o[17]) );
  LATCHX1_LVT \pc_o_reg[16]  ( .CLK(n40), .D(N35), .Q(pc_o[16]) );
  LATCHX1_LVT \pc_o_reg[15]  ( .CLK(n40), .D(N34), .Q(pc_o[15]) );
  LATCHX1_LVT \pc_o_reg[14]  ( .CLK(n40), .D(N33), .Q(pc_o[14]) );
  LATCHX1_LVT \pc_o_reg[13]  ( .CLK(n40), .D(N32), .Q(pc_o[13]) );
  LATCHX1_LVT \pc_o_reg[12]  ( .CLK(n40), .D(N31), .Q(pc_o[12]) );
  LATCHX1_LVT \pc_o_reg[11]  ( .CLK(n40), .D(N30), .Q(pc_o[11]) );
  LATCHX1_LVT \pc_o_reg[10]  ( .CLK(n40), .D(N29), .Q(pc_o[10]) );
  LATCHX1_LVT \pc_o_reg[9]  ( .CLK(n40), .D(N28), .Q(pc_o[9]) );
  LATCHX1_LVT \pc_o_reg[8]  ( .CLK(n40), .D(N27), .Q(pc_o[8]) );
  LATCHX1_LVT \pc_o_reg[7]  ( .CLK(n40), .D(N26), .Q(pc_o[7]) );
  LATCHX1_LVT \pc_o_reg[6]  ( .CLK(n40), .D(N25), .Q(pc_o[6]) );
  LATCHX1_LVT \pc_o_reg[5]  ( .CLK(n40), .D(N24), .Q(pc_o[5]) );
  LATCHX1_LVT \pc_o_reg[4]  ( .CLK(n40), .D(N23), .Q(pc_o[4]) );
  LATCHX1_LVT \pc_o_reg[3]  ( .CLK(n40), .D(N22), .Q(pc_o[3]) );
  LATCHX1_LVT \pc_o_reg[2]  ( .CLK(n40), .D(N21), .Q(pc_o[2]) );
  LATCHX1_LVT \pc_o_reg[1]  ( .CLK(n40), .D(N20), .Q(pc_o[1]) );
  LATCHX1_LVT mem_taking_reg ( .CLK(N16), .D(n43), .Q(mem_taking) );
  LATCHX1_LVT mem_re_reg ( .CLK(n6), .D(n43), .Q(mem_re) );
  LATCHX1_LVT stallreq_reg ( .CLK(N14), .D(N15), .Q(stallreq) );
  LATCHX1_LVT \mem_addr_o_reg[31]  ( .CLK(n42), .D(N116), .Q(mem_addr_o[31])
         );
  LATCHX1_LVT \mem_addr_o_reg[30]  ( .CLK(n42), .D(N115), .Q(mem_addr_o[30])
         );
  LATCHX1_LVT \mem_addr_o_reg[29]  ( .CLK(n42), .D(N114), .Q(mem_addr_o[29])
         );
  LATCHX1_LVT \mem_addr_o_reg[28]  ( .CLK(n42), .D(N113), .Q(mem_addr_o[28])
         );
  LATCHX1_LVT \mem_addr_o_reg[27]  ( .CLK(n6), .D(N112), .Q(mem_addr_o[27]) );
  LATCHX1_LVT \mem_addr_o_reg[26]  ( .CLK(n42), .D(N111), .Q(mem_addr_o[26])
         );
  LATCHX1_LVT \mem_addr_o_reg[25]  ( .CLK(n42), .D(N110), .Q(mem_addr_o[25])
         );
  LATCHX1_LVT \mem_addr_o_reg[24]  ( .CLK(n42), .D(N109), .Q(mem_addr_o[24])
         );
  LATCHX1_LVT \mem_addr_o_reg[23]  ( .CLK(n6), .D(N108), .Q(mem_addr_o[23]) );
  LATCHX1_LVT \mem_addr_o_reg[22]  ( .CLK(n6), .D(N107), .Q(mem_addr_o[22]) );
  LATCHX1_LVT \mem_addr_o_reg[21]  ( .CLK(n42), .D(N106), .Q(mem_addr_o[21])
         );
  LATCHX1_LVT \mem_addr_o_reg[20]  ( .CLK(n42), .D(N105), .Q(mem_addr_o[20])
         );
  LATCHX1_LVT \mem_addr_o_reg[19]  ( .CLK(n42), .D(N104), .Q(mem_addr_o[19])
         );
  LATCHX1_LVT \mem_addr_o_reg[18]  ( .CLK(n6), .D(N103), .Q(mem_addr_o[18]) );
  LATCHX1_LVT \mem_addr_o_reg[17]  ( .CLK(n6), .D(N102), .Q(mem_addr_o[17]) );
  LATCHX1_LVT \mem_addr_o_reg[16]  ( .CLK(n6), .D(N101), .Q(mem_addr_o[16]) );
  LATCHX1_LVT \mem_addr_o_reg[15]  ( .CLK(n6), .D(N100), .Q(mem_addr_o[15]) );
  LATCHX1_LVT \mem_addr_o_reg[14]  ( .CLK(n6), .D(N99), .Q(mem_addr_o[14]) );
  LATCHX1_LVT \mem_addr_o_reg[13]  ( .CLK(n6), .D(N98), .Q(mem_addr_o[13]) );
  LATCHX1_LVT \mem_addr_o_reg[12]  ( .CLK(n6), .D(N97), .Q(mem_addr_o[12]) );
  LATCHX1_LVT \mem_addr_o_reg[11]  ( .CLK(n6), .D(N96), .Q(mem_addr_o[11]) );
  LATCHX1_LVT \mem_addr_o_reg[10]  ( .CLK(n6), .D(N95), .Q(mem_addr_o[10]) );
  LATCHX1_LVT \mem_addr_o_reg[9]  ( .CLK(n6), .D(N94), .Q(mem_addr_o[9]) );
  LATCHX1_LVT \mem_addr_o_reg[8]  ( .CLK(n6), .D(N93), .Q(mem_addr_o[8]) );
  LATCHX1_LVT \mem_addr_o_reg[7]  ( .CLK(n6), .D(N92), .Q(mem_addr_o[7]) );
  LATCHX1_LVT \mem_addr_o_reg[6]  ( .CLK(n6), .D(N91), .Q(mem_addr_o[6]) );
  LATCHX1_LVT \mem_addr_o_reg[5]  ( .CLK(n6), .D(N90), .Q(mem_addr_o[5]) );
  LATCHX1_LVT \mem_addr_o_reg[4]  ( .CLK(n6), .D(N89), .Q(mem_addr_o[4]) );
  LATCHX1_LVT \mem_addr_o_reg[3]  ( .CLK(n6), .D(N88), .Q(mem_addr_o[3]) );
  LATCHX1_LVT \mem_addr_o_reg[2]  ( .CLK(n6), .D(N87), .Q(mem_addr_o[2]) );
  LATCHX1_LVT \mem_addr_o_reg[1]  ( .CLK(n6), .D(N86), .Q(mem_addr_o[1]) );
  LATCHX1_LVT \mem_addr_o_reg[0]  ( .CLK(n6), .D(N85), .Q(mem_addr_o[0]) );
  OR3X1_LVT U3 ( .A1(rst), .A2(br), .A3(right_one), .Y(N118) );
  INVX1_LVT U6 ( .A(right_one), .Y(n1) );
  NAND2X0_LVT U7 ( .A1(waiting_one), .A2(n1), .Y(n2) );
  NAND3X0_LVT U8 ( .A1(n36), .A2(n35), .A3(n2), .Y(n12) );
  NOR4X1_LVT U9 ( .A1(mem_busy[0]), .A2(mem_taking), .A3(mem_busy[1]), .A4(n12), .Y(n5) );
  INVX1_LVT U15 ( .A(mem_taking), .Y(n13) );
  NOR4X1_LVT U16 ( .A1(mem_busy[0]), .A2(mem_busy[1]), .A3(n13), .A4(n12), .Y(
        n15) );
  OR3X1_LVT U19 ( .A1(rst), .A2(br), .A3(n38), .Y(n9) );
  INVX1_LVT U29 ( .A(n12), .Y(n14) );
  AO222X1_LVT U30 ( .A1(n14), .A2(mem_busy[0]), .A3(n14), .A4(mem_busy[1]), 
        .A5(n14), .A6(n13), .Y(N15) );
  AND2X1_LVT U33 ( .A1(n37), .A2(mem_data_i[0]), .Y(N51) );
  AND2X1_LVT U34 ( .A1(n37), .A2(mem_data_i[1]), .Y(N52) );
  AND2X1_LVT U35 ( .A1(n37), .A2(mem_data_i[2]), .Y(N53) );
  AND2X1_LVT U36 ( .A1(n37), .A2(mem_data_i[3]), .Y(N54) );
  AND2X1_LVT U37 ( .A1(n37), .A2(mem_data_i[4]), .Y(N55) );
  AND2X1_LVT U38 ( .A1(n37), .A2(mem_data_i[5]), .Y(N56) );
  AND2X1_LVT U39 ( .A1(n37), .A2(mem_data_i[6]), .Y(N57) );
  AND2X1_LVT U40 ( .A1(n37), .A2(mem_data_i[7]), .Y(N58) );
  AND2X1_LVT U41 ( .A1(n37), .A2(mem_data_i[8]), .Y(N59) );
  AND2X1_LVT U42 ( .A1(n37), .A2(mem_data_i[9]), .Y(N60) );
  AND2X1_LVT U43 ( .A1(n37), .A2(mem_data_i[10]), .Y(N61) );
  AND2X1_LVT U44 ( .A1(n37), .A2(mem_data_i[11]), .Y(N62) );
  AND2X1_LVT U45 ( .A1(n37), .A2(mem_data_i[12]), .Y(N63) );
  AND2X1_LVT U46 ( .A1(n37), .A2(mem_data_i[13]), .Y(N64) );
  AND2X1_LVT U47 ( .A1(n37), .A2(mem_data_i[14]), .Y(N65) );
  AND2X1_LVT U49 ( .A1(n37), .A2(mem_data_i[15]), .Y(N66) );
  AND2X1_LVT U50 ( .A1(n37), .A2(mem_data_i[16]), .Y(N67) );
  AND2X1_LVT U51 ( .A1(n37), .A2(mem_data_i[17]), .Y(N68) );
  AND2X1_LVT U52 ( .A1(n37), .A2(mem_data_i[18]), .Y(N69) );
  AND2X1_LVT U53 ( .A1(n37), .A2(mem_data_i[19]), .Y(N70) );
  AND2X1_LVT U54 ( .A1(n37), .A2(mem_data_i[20]), .Y(N71) );
  AND2X1_LVT U55 ( .A1(n37), .A2(mem_data_i[21]), .Y(N72) );
  AND2X1_LVT U56 ( .A1(n37), .A2(mem_data_i[22]), .Y(N73) );
  AND2X1_LVT U57 ( .A1(n37), .A2(mem_data_i[23]), .Y(N74) );
  AND2X1_LVT U58 ( .A1(n37), .A2(mem_data_i[24]), .Y(N75) );
  AND2X1_LVT U59 ( .A1(n37), .A2(mem_data_i[25]), .Y(N76) );
  AND2X1_LVT U60 ( .A1(n37), .A2(mem_data_i[26]), .Y(N77) );
  AND2X1_LVT U61 ( .A1(n37), .A2(mem_data_i[27]), .Y(N78) );
  AND2X1_LVT U62 ( .A1(n37), .A2(mem_data_i[28]), .Y(N79) );
  AND2X1_LVT U63 ( .A1(n37), .A2(mem_data_i[29]), .Y(N80) );
  AND2X1_LVT U64 ( .A1(n37), .A2(mem_data_i[30]), .Y(N81) );
  AND2X1_LVT U65 ( .A1(n37), .A2(mem_data_i[31]), .Y(N82) );
  AND2X1_LVT U67 ( .A1(n38), .A2(pc_i[0]), .Y(N19) );
  AND2X1_LVT U68 ( .A1(n38), .A2(pc_i[1]), .Y(N20) );
  AND2X1_LVT U69 ( .A1(n38), .A2(pc_i[2]), .Y(N21) );
  AND2X1_LVT U70 ( .A1(n38), .A2(pc_i[3]), .Y(N22) );
  AND2X1_LVT U71 ( .A1(n38), .A2(pc_i[4]), .Y(N23) );
  AND2X1_LVT U72 ( .A1(n38), .A2(pc_i[5]), .Y(N24) );
  AND2X1_LVT U73 ( .A1(n38), .A2(pc_i[6]), .Y(N25) );
  AND2X1_LVT U74 ( .A1(n38), .A2(pc_i[7]), .Y(N26) );
  AND2X1_LVT U75 ( .A1(n38), .A2(pc_i[8]), .Y(N27) );
  AND2X1_LVT U76 ( .A1(n38), .A2(pc_i[9]), .Y(N28) );
  AND2X1_LVT U77 ( .A1(n38), .A2(pc_i[10]), .Y(N29) );
  AND2X1_LVT U78 ( .A1(n38), .A2(pc_i[11]), .Y(N30) );
  AND2X1_LVT U79 ( .A1(n38), .A2(pc_i[12]), .Y(N31) );
  AND2X1_LVT U80 ( .A1(n38), .A2(pc_i[13]), .Y(N32) );
  AND2X1_LVT U81 ( .A1(n38), .A2(pc_i[14]), .Y(N33) );
  AND2X1_LVT U82 ( .A1(n38), .A2(pc_i[15]), .Y(N34) );
  AND2X1_LVT U83 ( .A1(n38), .A2(pc_i[16]), .Y(N35) );
  AND2X1_LVT U84 ( .A1(n38), .A2(pc_i[17]), .Y(N36) );
  AND2X1_LVT U85 ( .A1(n38), .A2(pc_i[18]), .Y(N37) );
  AND2X1_LVT U86 ( .A1(n38), .A2(pc_i[19]), .Y(N38) );
  AND2X1_LVT U87 ( .A1(n38), .A2(pc_i[20]), .Y(N39) );
  AND2X1_LVT U88 ( .A1(n38), .A2(pc_i[21]), .Y(N40) );
  AND2X1_LVT U89 ( .A1(n38), .A2(pc_i[22]), .Y(N41) );
  AND2X1_LVT U90 ( .A1(n38), .A2(pc_i[23]), .Y(N42) );
  AND2X1_LVT U91 ( .A1(n38), .A2(pc_i[24]), .Y(N43) );
  AND2X1_LVT U92 ( .A1(n38), .A2(pc_i[25]), .Y(N44) );
  AND2X1_LVT U93 ( .A1(n38), .A2(pc_i[26]), .Y(N45) );
  AND2X1_LVT U94 ( .A1(n38), .A2(pc_i[27]), .Y(N46) );
  AND2X1_LVT U95 ( .A1(n38), .A2(pc_i[28]), .Y(N47) );
  AND2X1_LVT U96 ( .A1(n38), .A2(pc_i[29]), .Y(N48) );
  AND2X1_LVT U97 ( .A1(n38), .A2(pc_i[30]), .Y(N49) );
  AND2X1_LVT U98 ( .A1(n38), .A2(pc_i[31]), .Y(N50) );
  AND2X1_LVT U99 ( .A1(n43), .A2(pc_i[0]), .Y(N85) );
  AND2X1_LVT U101 ( .A1(n43), .A2(pc_i[1]), .Y(N86) );
  AND2X1_LVT U102 ( .A1(n43), .A2(pc_i[2]), .Y(N87) );
  AND2X1_LVT U104 ( .A1(n43), .A2(pc_i[3]), .Y(N88) );
  AND2X1_LVT U105 ( .A1(n43), .A2(pc_i[4]), .Y(N89) );
  AND2X1_LVT U106 ( .A1(n43), .A2(pc_i[5]), .Y(N90) );
  AND2X1_LVT U107 ( .A1(n43), .A2(pc_i[6]), .Y(N91) );
  AND2X1_LVT U108 ( .A1(n41), .A2(pc_i[7]), .Y(N92) );
  AND2X1_LVT U109 ( .A1(n5), .A2(pc_i[8]), .Y(N93) );
  AND2X1_LVT U110 ( .A1(n43), .A2(pc_i[9]), .Y(N94) );
  AND2X1_LVT U111 ( .A1(n43), .A2(pc_i[10]), .Y(N95) );
  AND2X1_LVT U112 ( .A1(n43), .A2(pc_i[11]), .Y(N96) );
  AND2X1_LVT U113 ( .A1(n43), .A2(pc_i[12]), .Y(N97) );
  AND2X1_LVT U114 ( .A1(n43), .A2(pc_i[13]), .Y(N98) );
  AND2X1_LVT U115 ( .A1(n43), .A2(pc_i[14]), .Y(N99) );
  AND2X1_LVT U116 ( .A1(n43), .A2(pc_i[15]), .Y(N100) );
  AND2X1_LVT U117 ( .A1(n43), .A2(pc_i[16]), .Y(N101) );
  AND2X1_LVT U118 ( .A1(n43), .A2(pc_i[17]), .Y(N102) );
  AND2X1_LVT U119 ( .A1(n43), .A2(pc_i[18]), .Y(N103) );
  AND2X1_LVT U120 ( .A1(n43), .A2(pc_i[19]), .Y(N104) );
  AND2X1_LVT U121 ( .A1(n43), .A2(pc_i[20]), .Y(N105) );
  AND2X1_LVT U122 ( .A1(n43), .A2(pc_i[21]), .Y(N106) );
  AND2X1_LVT U123 ( .A1(n43), .A2(pc_i[22]), .Y(N107) );
  AND2X1_LVT U124 ( .A1(n43), .A2(pc_i[23]), .Y(N108) );
  AND2X1_LVT U125 ( .A1(n43), .A2(pc_i[24]), .Y(N109) );
  AND2X1_LVT U126 ( .A1(n43), .A2(pc_i[25]), .Y(N110) );
  AND2X1_LVT U127 ( .A1(n43), .A2(pc_i[26]), .Y(N111) );
  AND2X1_LVT U128 ( .A1(n43), .A2(pc_i[27]), .Y(N112) );
  AND2X1_LVT U129 ( .A1(n43), .A2(pc_i[28]), .Y(N113) );
  AND2X1_LVT U130 ( .A1(n43), .A2(pc_i[29]), .Y(N114) );
  AND2X1_LVT U131 ( .A1(n43), .A2(pc_i[30]), .Y(N115) );
  AND2X1_LVT U132 ( .A1(n43), .A2(pc_i[31]), .Y(N116) );
  OR2X1_LVT U133 ( .A1(n40), .A2(n43), .Y(N16) );
  INVX1_LVT U134 ( .A(N118), .Y(n24) );
  NAND2X0_LVT U135 ( .A1(waiting_one), .A2(n24), .Y(N14) );
  AND2X1_LVT U137 ( .A1(br), .A2(n35), .Y(N119) );
  INVX1_LVT U4 ( .A(rst), .Y(n35) );
  INVX1_LVT U5 ( .A(br), .Y(n36) );
  NBUFFX8_LVT U10 ( .A(n15), .Y(n37) );
  NBUFFX8_LVT U11 ( .A(n15), .Y(n38) );
  NBUFFX8_LVT U13 ( .A(n9), .Y(n39) );
  NBUFFX8_LVT U14 ( .A(n9), .Y(n40) );
  OR2X4_LVT U12 ( .A1(rst), .A2(n43), .Y(n6) );
  NBUFFX4_LVT U17 ( .A(n5), .Y(n41) );
  NBUFFX4_LVT U18 ( .A(n6), .Y(n42) );
  NBUFFX4_LVT U20 ( .A(n41), .Y(n43) );
endmodule


module pipe_if_id ( clk, rst, if_pc, if_inst, stall, br, id_pc, id_inst );
  input [31:0] if_pc;
  input [31:0] if_inst;
  input [5:0] stall;
  output [31:0] id_pc;
  output [31:0] id_inst;
  input clk, rst, br;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n1, n72, n73, n82, n83, n84, n85;

  DFFX1_LVT \id_pc_reg[31]  ( .D(n35), .CLK(clk), .Q(id_pc[31]) );
  DFFX1_LVT \id_pc_reg[28]  ( .D(n32), .CLK(clk), .Q(id_pc[28]) );
  DFFX1_LVT \id_pc_reg[26]  ( .D(n30), .CLK(clk), .Q(id_pc[26]) );
  DFFX1_LVT \id_pc_reg[23]  ( .D(n27), .CLK(clk), .Q(id_pc[23]) );
  DFFX1_LVT \id_pc_reg[3]  ( .D(n7), .CLK(clk), .Q(id_pc[3]) );
  DFFX1_LVT \id_pc_reg[2]  ( .D(n6), .CLK(clk), .Q(id_pc[2]) );
  DFFX1_LVT \id_inst_reg[15]  ( .D(n51), .CLK(clk), .Q(id_inst[15]) );
  DFFX1_LVT \id_inst_reg[16]  ( .D(n52), .CLK(clk), .Q(id_inst[16]) );
  DFFX1_LVT \id_inst_reg[18]  ( .D(n54), .CLK(clk), .Q(id_inst[18]) );
  DFFX1_LVT \id_inst_reg[17]  ( .D(n53), .CLK(clk), .Q(id_inst[17]) );
  DFFX1_LVT \id_inst_reg[19]  ( .D(n55), .CLK(clk), .Q(id_inst[19]) );
  DFFX1_LVT \id_inst_reg[26]  ( .D(n62), .CLK(clk), .Q(id_inst[26]) );
  DFFX1_LVT \id_inst_reg[27]  ( .D(n63), .CLK(clk), .Q(id_inst[27]) );
  DFFX1_LVT \id_inst_reg[13]  ( .D(n49), .CLK(clk), .Q(id_inst[13]) );
  DFFX1_LVT \id_inst_reg[5]  ( .D(n41), .CLK(clk), .Q(id_inst[5]) );
  DFFX1_LVT \id_inst_reg[25]  ( .D(n61), .CLK(clk), .Q(id_inst[25]) );
  DFFX1_LVT \id_inst_reg[29]  ( .D(n65), .CLK(clk), .Q(id_inst[29]) );
  DFFX1_LVT \id_inst_reg[31]  ( .D(n67), .CLK(clk), .Q(id_inst[31]) );
  DFFX1_LVT \id_inst_reg[28]  ( .D(n64), .CLK(clk), .Q(id_inst[28]) );
  DFFX1_LVT \id_inst_reg[6]  ( .D(n42), .CLK(clk), .Q(id_inst[6]) );
  DFFX1_LVT \id_inst_reg[0]  ( .D(n36), .CLK(clk), .Q(id_inst[0]) );
  DFFX1_LVT \id_inst_reg[1]  ( .D(n37), .CLK(clk), .Q(id_inst[1]) );
  DFFX1_LVT \id_inst_reg[4]  ( .D(n40), .CLK(clk), .Q(id_inst[4]) );
  DFFX1_LVT \id_inst_reg[2]  ( .D(n38), .CLK(clk), .Q(id_inst[2]) );
  DFFX1_LVT \id_inst_reg[3]  ( .D(n39), .CLK(clk), .Q(id_inst[3]) );
  NOR3X0_LVT U3 ( .A1(stall[1]), .A2(rst), .A3(br), .Y(n72) );
  NOR2X0_LVT U6 ( .A1(rst), .A2(br), .Y(n1) );
  AND3X1_LVT U7 ( .A1(stall[1]), .A2(n1), .A3(stall[2]), .Y(n73) );
  AO22X1_LVT U10 ( .A1(n84), .A2(if_inst[31]), .A3(n82), .A4(id_inst[31]), .Y(
        n67) );
  AO22X1_LVT U11 ( .A1(n84), .A2(if_inst[30]), .A3(n82), .A4(id_inst[30]), .Y(
        n66) );
  AO22X1_LVT U12 ( .A1(n84), .A2(if_inst[29]), .A3(n82), .A4(id_inst[29]), .Y(
        n65) );
  AO22X1_LVT U13 ( .A1(n84), .A2(if_inst[28]), .A3(n82), .A4(id_inst[28]), .Y(
        n64) );
  AO22X1_LVT U14 ( .A1(n84), .A2(if_inst[27]), .A3(n82), .A4(id_inst[27]), .Y(
        n63) );
  AO22X1_LVT U15 ( .A1(n84), .A2(if_inst[26]), .A3(n82), .A4(id_inst[26]), .Y(
        n62) );
  AO22X1_LVT U16 ( .A1(n84), .A2(if_inst[25]), .A3(n82), .A4(id_inst[25]), .Y(
        n61) );
  AO22X1_LVT U17 ( .A1(n84), .A2(if_inst[24]), .A3(n82), .A4(id_inst[24]), .Y(
        n60) );
  AO22X1_LVT U18 ( .A1(n84), .A2(if_inst[23]), .A3(n82), .A4(id_inst[23]), .Y(
        n59) );
  AO22X1_LVT U19 ( .A1(n84), .A2(if_inst[22]), .A3(n82), .A4(id_inst[22]), .Y(
        n58) );
  AO22X1_LVT U20 ( .A1(n84), .A2(if_inst[21]), .A3(n82), .A4(id_inst[21]), .Y(
        n57) );
  AO22X1_LVT U21 ( .A1(n84), .A2(if_inst[20]), .A3(n82), .A4(id_inst[20]), .Y(
        n56) );
  AO22X1_LVT U22 ( .A1(n84), .A2(if_inst[19]), .A3(n82), .A4(id_inst[19]), .Y(
        n55) );
  AO22X1_LVT U23 ( .A1(n84), .A2(if_inst[18]), .A3(n82), .A4(id_inst[18]), .Y(
        n54) );
  AO22X1_LVT U24 ( .A1(n84), .A2(if_inst[17]), .A3(n82), .A4(id_inst[17]), .Y(
        n53) );
  AO22X1_LVT U27 ( .A1(n84), .A2(if_inst[16]), .A3(n82), .A4(id_inst[16]), .Y(
        n52) );
  AO22X1_LVT U28 ( .A1(n84), .A2(if_inst[15]), .A3(n82), .A4(id_inst[15]), .Y(
        n51) );
  AO22X1_LVT U29 ( .A1(n84), .A2(if_inst[14]), .A3(n82), .A4(id_inst[14]), .Y(
        n50) );
  AO22X1_LVT U30 ( .A1(n84), .A2(if_inst[13]), .A3(n82), .A4(id_inst[13]), .Y(
        n49) );
  AO22X1_LVT U31 ( .A1(n84), .A2(if_inst[12]), .A3(n82), .A4(id_inst[12]), .Y(
        n48) );
  AO22X1_LVT U32 ( .A1(n84), .A2(if_inst[11]), .A3(n82), .A4(id_inst[11]), .Y(
        n47) );
  AO22X1_LVT U33 ( .A1(n84), .A2(if_inst[10]), .A3(n82), .A4(id_inst[10]), .Y(
        n46) );
  AO22X1_LVT U34 ( .A1(n84), .A2(if_inst[9]), .A3(n82), .A4(id_inst[9]), .Y(
        n45) );
  AO22X1_LVT U35 ( .A1(n84), .A2(if_inst[8]), .A3(n82), .A4(id_inst[8]), .Y(
        n44) );
  AO22X1_LVT U36 ( .A1(n84), .A2(if_inst[7]), .A3(n82), .A4(id_inst[7]), .Y(
        n43) );
  AO22X1_LVT U37 ( .A1(n84), .A2(if_inst[6]), .A3(n82), .A4(id_inst[6]), .Y(
        n42) );
  AO22X1_LVT U38 ( .A1(n84), .A2(if_inst[5]), .A3(n82), .A4(id_inst[5]), .Y(
        n41) );
  AO22X1_LVT U39 ( .A1(n84), .A2(if_inst[4]), .A3(n82), .A4(id_inst[4]), .Y(
        n40) );
  AO22X1_LVT U40 ( .A1(n84), .A2(if_inst[3]), .A3(n82), .A4(id_inst[3]), .Y(
        n39) );
  AO22X1_LVT U41 ( .A1(n84), .A2(if_inst[2]), .A3(n82), .A4(id_inst[2]), .Y(
        n38) );
  AO22X1_LVT U46 ( .A1(n84), .A2(if_inst[1]), .A3(n82), .A4(id_inst[1]), .Y(
        n37) );
  AO22X1_LVT U47 ( .A1(n84), .A2(if_inst[0]), .A3(n82), .A4(id_inst[0]), .Y(
        n36) );
  AO22X1_LVT U48 ( .A1(n85), .A2(if_pc[31]), .A3(n83), .A4(id_pc[31]), .Y(n35)
         );
  AO22X1_LVT U49 ( .A1(n85), .A2(if_pc[30]), .A3(n83), .A4(id_pc[30]), .Y(n34)
         );
  AO22X1_LVT U50 ( .A1(n85), .A2(if_pc[29]), .A3(n83), .A4(id_pc[29]), .Y(n33)
         );
  AO22X1_LVT U51 ( .A1(n85), .A2(if_pc[28]), .A3(n83), .A4(id_pc[28]), .Y(n32)
         );
  AO22X1_LVT U52 ( .A1(n85), .A2(if_pc[27]), .A3(n83), .A4(id_pc[27]), .Y(n31)
         );
  AO22X1_LVT U53 ( .A1(n85), .A2(if_pc[26]), .A3(n83), .A4(id_pc[26]), .Y(n30)
         );
  AO22X1_LVT U54 ( .A1(n85), .A2(if_pc[25]), .A3(n83), .A4(id_pc[25]), .Y(n29)
         );
  AO22X1_LVT U55 ( .A1(n85), .A2(if_pc[24]), .A3(n83), .A4(id_pc[24]), .Y(n28)
         );
  AO22X1_LVT U56 ( .A1(n85), .A2(if_pc[23]), .A3(n83), .A4(id_pc[23]), .Y(n27)
         );
  AO22X1_LVT U57 ( .A1(n85), .A2(if_pc[22]), .A3(n83), .A4(id_pc[22]), .Y(n26)
         );
  AO22X1_LVT U58 ( .A1(n85), .A2(if_pc[21]), .A3(n83), .A4(id_pc[21]), .Y(n25)
         );
  AO22X1_LVT U59 ( .A1(n85), .A2(if_pc[20]), .A3(n83), .A4(id_pc[20]), .Y(n24)
         );
  AO22X1_LVT U60 ( .A1(n85), .A2(if_pc[19]), .A3(n83), .A4(id_pc[19]), .Y(n23)
         );
  AO22X1_LVT U63 ( .A1(n85), .A2(if_pc[18]), .A3(n83), .A4(id_pc[18]), .Y(n22)
         );
  AO22X1_LVT U64 ( .A1(n85), .A2(if_pc[17]), .A3(n83), .A4(id_pc[17]), .Y(n21)
         );
  AO22X1_LVT U65 ( .A1(n85), .A2(if_pc[16]), .A3(n83), .A4(id_pc[16]), .Y(n20)
         );
  AO22X1_LVT U66 ( .A1(n85), .A2(if_pc[15]), .A3(n83), .A4(id_pc[15]), .Y(n19)
         );
  AO22X1_LVT U67 ( .A1(n85), .A2(if_pc[14]), .A3(n83), .A4(id_pc[14]), .Y(n18)
         );
  AO22X1_LVT U68 ( .A1(n85), .A2(if_pc[13]), .A3(n83), .A4(id_pc[13]), .Y(n17)
         );
  AO22X1_LVT U69 ( .A1(n85), .A2(if_pc[12]), .A3(n83), .A4(id_pc[12]), .Y(n16)
         );
  AO22X1_LVT U70 ( .A1(n85), .A2(if_pc[11]), .A3(n83), .A4(id_pc[11]), .Y(n15)
         );
  AO22X1_LVT U71 ( .A1(n85), .A2(if_pc[10]), .A3(n83), .A4(id_pc[10]), .Y(n14)
         );
  AO22X1_LVT U72 ( .A1(n85), .A2(if_pc[9]), .A3(n83), .A4(id_pc[9]), .Y(n13)
         );
  AO22X1_LVT U73 ( .A1(n85), .A2(if_pc[8]), .A3(n83), .A4(id_pc[8]), .Y(n12)
         );
  AO22X1_LVT U74 ( .A1(n85), .A2(if_pc[7]), .A3(n83), .A4(id_pc[7]), .Y(n11)
         );
  AO22X1_LVT U75 ( .A1(n85), .A2(if_pc[6]), .A3(n83), .A4(id_pc[6]), .Y(n10)
         );
  AO22X1_LVT U76 ( .A1(n85), .A2(if_pc[5]), .A3(n83), .A4(id_pc[5]), .Y(n9) );
  AO22X1_LVT U77 ( .A1(n85), .A2(if_pc[4]), .A3(n83), .A4(id_pc[4]), .Y(n8) );
  AO22X1_LVT U80 ( .A1(n85), .A2(if_pc[3]), .A3(n83), .A4(id_pc[3]), .Y(n7) );
  AO22X1_LVT U81 ( .A1(n85), .A2(if_pc[2]), .A3(n83), .A4(id_pc[2]), .Y(n6) );
  AO22X1_LVT U82 ( .A1(n85), .A2(if_pc[1]), .A3(n83), .A4(id_pc[1]), .Y(n5) );
  AO22X1_LVT U83 ( .A1(n85), .A2(if_pc[0]), .A3(n83), .A4(id_pc[0]), .Y(n4) );
  NBUFFX8_LVT U4 ( .A(n73), .Y(n82) );
  NBUFFX8_LVT U5 ( .A(n73), .Y(n83) );
  NBUFFX8_LVT U8 ( .A(n72), .Y(n84) );
  NBUFFX8_LVT U9 ( .A(n72), .Y(n85) );
  DFFX2_LVT \id_pc_reg[10]  ( .D(n14), .CLK(clk), .Q(id_pc[10]) );
  DFFX2_LVT \id_pc_reg[11]  ( .D(n15), .CLK(clk), .Q(id_pc[11]) );
  DFFX2_LVT \id_pc_reg[14]  ( .D(n18), .CLK(clk), .Q(id_pc[14]) );
  DFFX2_LVT \id_pc_reg[12]  ( .D(n16), .CLK(clk), .Q(id_pc[12]) );
  DFFX2_LVT \id_pc_reg[13]  ( .D(n17), .CLK(clk), .Q(id_pc[13]) );
  DFFX2_LVT \id_pc_reg[6]  ( .D(n10), .CLK(clk), .Q(id_pc[6]) );
  DFFX2_LVT \id_pc_reg[7]  ( .D(n11), .CLK(clk), .Q(id_pc[7]) );
  DFFX2_LVT \id_pc_reg[9]  ( .D(n13), .CLK(clk), .Q(id_pc[9]) );
  DFFX2_LVT \id_inst_reg[24]  ( .D(n60), .CLK(clk), .Q(id_inst[24]) );
  DFFX2_LVT \id_pc_reg[8]  ( .D(n12), .CLK(clk), .Q(id_pc[8]) );
  DFFX2_LVT \id_pc_reg[16]  ( .D(n20), .CLK(clk), .Q(id_pc[16]) );
  DFFX2_LVT \id_pc_reg[4]  ( .D(n8), .CLK(clk), .Q(id_pc[4]) );
  DFFX2_LVT \id_pc_reg[5]  ( .D(n9), .CLK(clk), .Q(id_pc[5]) );
  DFFX2_LVT \id_inst_reg[21]  ( .D(n57), .CLK(clk), .Q(id_inst[21]) );
  DFFX2_LVT \id_inst_reg[30]  ( .D(n66), .CLK(clk), .Q(id_inst[30]) );
  DFFX2_LVT \id_pc_reg[17]  ( .D(n21), .CLK(clk), .Q(id_pc[17]) );
  DFFX2_LVT \id_pc_reg[15]  ( .D(n19), .CLK(clk), .Q(id_pc[15]) );
  DFFX2_LVT \id_pc_reg[18]  ( .D(n22), .CLK(clk), .Q(id_pc[18]) );
  DFFX2_LVT \id_inst_reg[22]  ( .D(n58), .CLK(clk), .Q(id_inst[22]) );
  DFFX2_LVT \id_inst_reg[20]  ( .D(n56), .CLK(clk), .Q(id_inst[20]) );
  DFFX2_LVT \id_inst_reg[23]  ( .D(n59), .CLK(clk), .Q(id_inst[23]) );
  DFFX2_LVT \id_pc_reg[20]  ( .D(n24), .CLK(clk), .Q(id_pc[20]) );
  DFFX2_LVT \id_pc_reg[19]  ( .D(n23), .CLK(clk), .Q(id_pc[19]) );
  DFFX2_LVT \id_pc_reg[21]  ( .D(n25), .CLK(clk), .Q(id_pc[21]) );
  DFFX2_LVT \id_pc_reg[22]  ( .D(n26), .CLK(clk), .Q(id_pc[22]) );
  DFFX2_LVT \id_inst_reg[12]  ( .D(n48), .CLK(clk), .Q(id_inst[12]) );
  DFFX2_LVT \id_pc_reg[30]  ( .D(n34), .CLK(clk), .Q(id_pc[30]) );
  DFFX2_LVT \id_pc_reg[24]  ( .D(n28), .CLK(clk), .Q(id_pc[24]) );
  DFFX2_LVT \id_pc_reg[29]  ( .D(n33), .CLK(clk), .Q(id_pc[29]) );
  DFFX2_LVT \id_inst_reg[14]  ( .D(n50), .CLK(clk), .Q(id_inst[14]) );
  DFFX2_LVT \id_pc_reg[25]  ( .D(n29), .CLK(clk), .Q(id_pc[25]) );
  DFFX2_LVT \id_pc_reg[1]  ( .D(n5), .CLK(clk), .Q(id_pc[1]) );
  DFFX2_LVT \id_pc_reg[27]  ( .D(n31), .CLK(clk), .Q(id_pc[27]) );
  DFFX2_LVT \id_pc_reg[0]  ( .D(n4), .CLK(clk), .Q(id_pc[0]) );
  DFFX2_LVT \id_inst_reg[7]  ( .D(n43), .CLK(clk), .Q(id_inst[7]) );
  DFFX2_LVT \id_inst_reg[10]  ( .D(n46), .CLK(clk), .Q(id_inst[10]) );
  DFFX2_LVT \id_inst_reg[9]  ( .D(n45), .CLK(clk), .Q(id_inst[9]) );
  DFFX2_LVT \id_inst_reg[8]  ( .D(n44), .CLK(clk), .Q(id_inst[8]) );
  DFFX2_LVT \id_inst_reg[11]  ( .D(n47), .CLK(clk), .Q(id_inst[11]) );
endmodule


module inst_decoder ( rst, pc, inst, reg_data1, reg_data2, ex_aluop, ex_we, 
        ex_reg_wdata, ex_reg_waddr, mem_we, mem_reg_wdata, mem_reg_waddr, re1, 
        re2, reg_addr1, reg_addr2, aluop, alusel, opv1, opv2, reg_waddr, we, 
        stallreq, br, br_addr, link_addr, mem_offset );
  input [31:0] pc;
  input [31:0] inst;
  input [31:0] reg_data1;
  input [31:0] reg_data2;
  input [7:0] ex_aluop;
  input [31:0] ex_reg_wdata;
  input [4:0] ex_reg_waddr;
  input [31:0] mem_reg_wdata;
  input [4:0] mem_reg_waddr;
  output [4:0] reg_addr1;
  output [4:0] reg_addr2;
  output [7:0] aluop;
  output [2:0] alusel;
  output [31:0] opv1;
  output [31:0] opv2;
  output [4:0] reg_waddr;
  output [31:0] br_addr;
  output [31:0] link_addr;
  output [31:0] mem_offset;
  input rst, ex_we, mem_we;
  output re1, re2, we, stallreq, br;
  wire   N94, N635, N636, N637, N638, N639, N640, N641, N642, N643, N644, N645,
         N646, N647, N648, N649, N650, N651, N652, N653, N654, N655, N656,
         N657, N658, N659, N660, N661, N662, N663, N664, N665, N666, N696,
         N697, N698, N699, N700, N701, N702, N703, N704, N705, N706, N707,
         N708, N709, N710, N711, N712, N713, N714, N715, N716, N717, N718,
         N719, N720, N721, N722, N723, N724, N725, N726, N727, n1, n2, n4, n5,
         n6, n7, n8, n10, n11, n12, n13, n14, n15, n16, n17, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n257, n258, n259, n260, n261, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n560,
         n561, n563, n565, n566, n568, n569, n570, n573, n574, n575, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n640, n641, n647, n648, n649, n650, n651, n653, n654, n655,
         n657, n658, n659, n661, n662, n663, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n703,
         n704, n705, n707, n708, n709, n712, n713, n714, n720, n721, n722,
         n723, n728, n730, n731, n732, n733, n734, n735, n736, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n754, n755, n756, n757, n758, n759, n760, n761, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n787, n788, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n829, n830, n831, n832,
         n833, n834, n835, n836, \mem_offset[11] , n838, n839;
  assign mem_offset[13] = mem_offset[31];
  assign mem_offset[14] = mem_offset[31];
  assign mem_offset[15] = mem_offset[31];
  assign mem_offset[16] = mem_offset[31];
  assign mem_offset[18] = mem_offset[31];
  assign mem_offset[21] = mem_offset[31];
  assign mem_offset[23] = mem_offset[31];
  assign mem_offset[24] = mem_offset[31];
  assign mem_offset[25] = mem_offset[31];
  assign mem_offset[28] = mem_offset[31];
  assign mem_offset[29] = mem_offset[31];
  assign mem_offset[30] = mem_offset[31];
  assign N94 = inst[14];
  assign mem_offset[27] = \mem_offset[11] ;
  assign mem_offset[20] = \mem_offset[11] ;
  assign mem_offset[17] = \mem_offset[11] ;
  assign mem_offset[22] = \mem_offset[11] ;
  assign mem_offset[19] = \mem_offset[11] ;
  assign mem_offset[12] = \mem_offset[11] ;
  assign mem_offset[26] = \mem_offset[11] ;
  assign mem_offset[11] = \mem_offset[11] ;

  LATCHX1_LVT \opv1_reg[31]  ( .CLK(n835), .D(N666), .Q(opv1[31]) );
  LATCHX1_LVT \opv1_reg[30]  ( .CLK(n237), .D(N665), .Q(opv1[30]) );
  LATCHX1_LVT \opv1_reg[29]  ( .CLK(n835), .D(N664), .Q(opv1[29]) );
  LATCHX1_LVT \opv1_reg[28]  ( .CLK(n237), .D(N663), .Q(opv1[28]) );
  LATCHX1_LVT \opv1_reg[27]  ( .CLK(n835), .D(N662), .Q(opv1[27]) );
  LATCHX1_LVT \opv1_reg[26]  ( .CLK(n835), .D(N661), .Q(opv1[26]) );
  LATCHX1_LVT \opv1_reg[24]  ( .CLK(n835), .D(N659), .Q(opv1[24]) );
  LATCHX1_LVT \opv1_reg[23]  ( .CLK(n835), .D(N658), .Q(opv1[23]) );
  LATCHX1_LVT \opv1_reg[22]  ( .CLK(n835), .D(N657), .Q(opv1[22]) );
  LATCHX1_LVT \opv1_reg[21]  ( .CLK(n835), .D(N656), .Q(opv1[21]) );
  LATCHX1_LVT \opv1_reg[20]  ( .CLK(n835), .D(N655), .Q(opv1[20]) );
  LATCHX1_LVT \opv1_reg[19]  ( .CLK(n835), .D(N654), .Q(opv1[19]) );
  LATCHX1_LVT \opv1_reg[18]  ( .CLK(n835), .D(N653), .Q(opv1[18]) );
  LATCHX1_LVT \opv1_reg[15]  ( .CLK(n835), .D(N650), .Q(opv1[15]) );
  LATCHX1_LVT \opv1_reg[14]  ( .CLK(n835), .D(N649), .Q(opv1[14]) );
  LATCHX1_LVT \opv1_reg[13]  ( .CLK(n835), .D(N648), .Q(opv1[13]) );
  LATCHX1_LVT \opv1_reg[12]  ( .CLK(n835), .D(N647), .Q(opv1[12]) );
  LATCHX1_LVT \opv1_reg[11]  ( .CLK(n835), .D(N646), .Q(opv1[11]) );
  LATCHX1_LVT \opv1_reg[10]  ( .CLK(n835), .D(N645), .Q(opv1[10]) );
  LATCHX1_LVT \opv1_reg[9]  ( .CLK(n835), .D(N644), .Q(opv1[9]) );
  LATCHX1_LVT \opv1_reg[8]  ( .CLK(n835), .D(N643), .Q(opv1[8]) );
  LATCHX1_LVT \opv1_reg[7]  ( .CLK(n835), .D(N642), .Q(opv1[7]) );
  LATCHX1_LVT \opv1_reg[6]  ( .CLK(n835), .D(N641), .Q(opv1[6]) );
  LATCHX1_LVT \opv1_reg[5]  ( .CLK(n835), .D(N640), .Q(opv1[5]) );
  LATCHX1_LVT \opv1_reg[4]  ( .CLK(n237), .D(N639), .Q(opv1[4]) );
  LATCHX1_LVT \opv1_reg[3]  ( .CLK(n237), .D(N638), .Q(opv1[3]) );
  LATCHX1_LVT \opv1_reg[2]  ( .CLK(n237), .D(N637), .Q(opv1[2]) );
  LATCHX1_LVT \opv1_reg[1]  ( .CLK(n237), .D(N636), .Q(opv1[1]) );
  LATCHX1_LVT \opv1_reg[0]  ( .CLK(n237), .D(N635), .Q(opv1[0]) );
  LATCHX1_LVT \opv2_reg[31]  ( .CLK(n254), .D(N727), .Q(opv2[31]) );
  LATCHX1_LVT \opv2_reg[30]  ( .CLK(n254), .D(N726), .Q(opv2[30]) );
  LATCHX1_LVT \opv2_reg[29]  ( .CLK(n254), .D(N725), .Q(opv2[29]) );
  LATCHX1_LVT \opv2_reg[28]  ( .CLK(n254), .D(N724), .Q(opv2[28]) );
  LATCHX1_LVT \opv2_reg[27]  ( .CLK(n838), .D(N723), .Q(opv2[27]) );
  LATCHX1_LVT \opv2_reg[26]  ( .CLK(n254), .D(N722), .Q(opv2[26]) );
  LATCHX1_LVT \opv2_reg[25]  ( .CLK(n838), .D(N721), .Q(opv2[25]) );
  LATCHX1_LVT \opv2_reg[24]  ( .CLK(n838), .D(N720), .Q(opv2[24]) );
  LATCHX1_LVT \opv2_reg[23]  ( .CLK(n838), .D(N719), .Q(opv2[23]) );
  LATCHX1_LVT \opv2_reg[22]  ( .CLK(n254), .D(N718), .Q(opv2[22]) );
  LATCHX1_LVT \opv2_reg[21]  ( .CLK(n838), .D(N717), .Q(opv2[21]) );
  LATCHX1_LVT \opv2_reg[20]  ( .CLK(n838), .D(N716), .Q(opv2[20]) );
  LATCHX1_LVT \opv2_reg[19]  ( .CLK(n838), .D(N715), .Q(opv2[19]) );
  LATCHX1_LVT \opv2_reg[18]  ( .CLK(n838), .D(N714), .Q(opv2[18]) );
  LATCHX1_LVT \opv2_reg[17]  ( .CLK(n838), .D(N713), .Q(opv2[17]) );
  LATCHX1_LVT \opv2_reg[16]  ( .CLK(n838), .D(N712), .Q(opv2[16]) );
  LATCHX1_LVT \opv2_reg[15]  ( .CLK(n254), .D(N711), .Q(opv2[15]) );
  LATCHX1_LVT \opv2_reg[14]  ( .CLK(n838), .D(N710), .Q(opv2[14]) );
  LATCHX1_LVT \opv2_reg[13]  ( .CLK(n838), .D(N709), .Q(opv2[13]) );
  LATCHX1_LVT \opv2_reg[12]  ( .CLK(n838), .D(N708), .Q(opv2[12]) );
  LATCHX1_LVT \opv2_reg[11]  ( .CLK(n838), .D(N707), .Q(opv2[11]) );
  LATCHX1_LVT \opv2_reg[10]  ( .CLK(n838), .D(N706), .Q(opv2[10]) );
  LATCHX1_LVT \opv2_reg[9]  ( .CLK(n838), .D(N705), .Q(opv2[9]) );
  LATCHX1_LVT \opv2_reg[8]  ( .CLK(n838), .D(N704), .Q(opv2[8]) );
  LATCHX1_LVT \opv2_reg[7]  ( .CLK(n838), .D(N703), .Q(opv2[7]) );
  LATCHX1_LVT \opv2_reg[6]  ( .CLK(n838), .D(N702), .Q(opv2[6]) );
  LATCHX1_LVT \opv2_reg[5]  ( .CLK(n838), .D(N701), .Q(opv2[5]) );
  LATCHX1_LVT \opv2_reg[4]  ( .CLK(n254), .D(N700), .Q(opv2[4]) );
  LATCHX1_LVT \opv2_reg[3]  ( .CLK(n254), .D(N699), .Q(opv2[3]) );
  LATCHX1_LVT \opv2_reg[2]  ( .CLK(n254), .D(N698), .Q(opv2[2]) );
  LATCHX1_LVT \opv2_reg[1]  ( .CLK(n254), .D(N697), .Q(opv2[1]) );
  LATCHX1_LVT \opv2_reg[0]  ( .CLK(n254), .D(N696), .Q(opv2[0]) );
  NAND3X0_LVT U4 ( .A1(inst[0]), .A2(inst[1]), .A3(n809), .Y(n756) );
  INVX1_LVT U5 ( .A(n756), .Y(n751) );
  INVX1_LVT U6 ( .A(inst[6]), .Y(n238) );
  AND3X1_LVT U8 ( .A1(n238), .A2(n811), .A3(inst[4]), .Y(n748) );
  INVX1_LVT U9 ( .A(inst[2]), .Y(n8) );
  NAND3X0_LVT U10 ( .A1(n751), .A2(n748), .A3(n8), .Y(n779) );
  INVX1_LVT U11 ( .A(n779), .Y(n765) );
  OR4X1_LVT U13 ( .A1(inst[28]), .A2(inst[31]), .A3(inst[29]), .A4(inst[25]), 
        .Y(n1) );
  OR3X1_LVT U14 ( .A1(inst[27]), .A2(inst[26]), .A3(n1), .Y(n758) );
  OA22X1_LVT U17 ( .A1(n812), .A2(n813), .A3(N94), .A4(inst[12]), .Y(n764) );
  INVX1_LVT U18 ( .A(n764), .Y(n760) );
  NAND3X0_LVT U19 ( .A1(n836), .A2(n758), .A3(n760), .Y(n2) );
  NAND3X0_LVT U20 ( .A1(inst[5]), .A2(n765), .A3(n2), .Y(n740) );
  NOR3X0_LVT U21 ( .A1(inst[3]), .A2(inst[2]), .A3(inst[4]), .Y(n492) );
  NAND4X0_LVT U22 ( .A1(n751), .A2(inst[6]), .A3(inst[5]), .A4(n492), .Y(n780)
         );
  INVX1_LVT U23 ( .A(n780), .Y(n802) );
  OR2X1_LVT U25 ( .A1(n814), .A2(N94), .Y(n744) );
  NAND2X0_LVT U26 ( .A1(n802), .A2(n744), .Y(n755) );
  AND4X1_LVT U27 ( .A1(inst[5]), .A2(n492), .A3(n238), .A4(n812), .Y(n754) );
  NAND2X0_LVT U28 ( .A1(inst[12]), .A2(inst[13]), .Y(n776) );
  AND2X1_LVT U29 ( .A1(n754), .A2(n776), .Y(n239) );
  NAND2X0_LVT U30 ( .A1(n751), .A2(n239), .Y(n799) );
  NAND3X0_LVT U31 ( .A1(n740), .A2(n755), .A3(n799), .Y(re2) );
  INVX1_LVT U32 ( .A(re2), .Y(n252) );
  NAND2X0_LVT U33 ( .A1(n252), .A2(n809), .Y(n243) );
  NAND2X0_LVT U34 ( .A1(inst[22]), .A2(n243), .Y(n260) );
  NAND2X0_LVT U36 ( .A1(inst[23]), .A2(n243), .Y(n246) );
  NAND2X0_LVT U38 ( .A1(inst[20]), .A2(n243), .Y(n248) );
  INVX1_LVT U39 ( .A(n248), .Y(reg_addr2[0]) );
  INVX1_LVT U40 ( .A(inst[5]), .Y(n269) );
  NAND4X0_LVT U41 ( .A1(n751), .A2(n492), .A3(n269), .A4(n238), .Y(n782) );
  INVX1_LVT U42 ( .A(n782), .Y(n796) );
  NAND2X0_LVT U43 ( .A1(n812), .A2(n813), .Y(n745) );
  NAND2X0_LVT U44 ( .A1(inst[13]), .A2(n745), .Y(n240) );
  NAND2X0_LVT U45 ( .A1(n796), .A2(n240), .Y(n731) );
  NAND4X0_LVT U46 ( .A1(inst[12]), .A2(N94), .A3(n836), .A4(n758), .Y(n4) );
  NAND3X0_LVT U47 ( .A1(n765), .A2(n269), .A3(n4), .Y(n309) );
  NAND2X0_LVT U48 ( .A1(n731), .A2(n309), .Y(n733) );
  INVX1_LVT U49 ( .A(n733), .Y(n13) );
  INVX1_LVT U50 ( .A(n243), .Y(n12) );
  AND2X1_LVT U51 ( .A1(inst[0]), .A2(inst[1]), .Y(n735) );
  INVX1_LVT U52 ( .A(inst[6]), .Y(n6) );
  INVX1_LVT U53 ( .A(inst[5]), .Y(n5) );
  OR2X1_LVT U54 ( .A1(n6), .A2(n5), .Y(n7) );
  NOR3X0_LVT U55 ( .A1(n8), .A2(inst[4]), .A3(n7), .Y(n746) );
  AND2X1_LVT U56 ( .A1(n746), .A2(n811), .Y(n10) );
  NAND2X0_LVT U59 ( .A1(n735), .A2(n823), .Y(n11) );
  NAND3X0_LVT U60 ( .A1(n13), .A2(n12), .A3(n11), .Y(n227) );
  NAND2X0_LVT U61 ( .A1(inst[16]), .A2(n227), .Y(n583) );
  INVX1_LVT U62 ( .A(n583), .Y(reg_addr1[1]) );
  NAND2X0_LVT U63 ( .A1(inst[19]), .A2(n227), .Y(n581) );
  NAND2X0_LVT U65 ( .A1(inst[18]), .A2(n227), .Y(n588) );
  INVX1_LVT U67 ( .A(n733), .Y(n16) );
  INVX1_LVT U68 ( .A(re2), .Y(n15) );
  NAND2X0_LVT U69 ( .A1(n751), .A2(n823), .Y(n14) );
  NAND3X0_LVT U70 ( .A1(n16), .A2(n15), .A3(n14), .Y(re1) );
  NAND2X0_LVT U71 ( .A1(inst[17]), .A2(n227), .Y(n582) );
  INVX1_LVT U74 ( .A(opv1[29]), .Y(n79) );
  INVX1_LVT U75 ( .A(opv1[28]), .Y(n78) );
  OR2X1_LVT U76 ( .A1(n78), .A2(opv2[28]), .Y(n182) );
  AO222X1_LVT U77 ( .A1(opv2[29]), .A2(n79), .A3(opv2[29]), .A4(n182), .A5(n79), .A6(n182), .Y(n85) );
  INVX1_LVT U78 ( .A(opv1[27]), .Y(n175) );
  INVX1_LVT U79 ( .A(opv1[26]), .Y(n73) );
  AOI22X1_LVT U80 ( .A1(n175), .A2(opv2[27]), .A3(n73), .A4(opv2[26]), .Y(n177) );
  NAND2X0_LVT U82 ( .A1(opv2[25]), .A2(n833), .Y(n17) );
  NAND2X0_LVT U83 ( .A1(n177), .A2(n17), .Y(n77) );
  OA22X1_LVT U85 ( .A1(opv2[25]), .A2(n833), .A3(opv2[24]), .A4(n832), .Y(n76)
         );
  INVX1_LVT U86 ( .A(n77), .Y(n21) );
  NAND2X0_LVT U87 ( .A1(opv2[24]), .A2(n832), .Y(n20) );
  NAND2X0_LVT U88 ( .A1(n21), .A2(n20), .Y(n198) );
  INVX1_LVT U89 ( .A(opv2[14]), .Y(n23) );
  INVX1_LVT U90 ( .A(opv2[15]), .Y(n102) );
  OA22X1_LVT U91 ( .A1(opv1[14]), .A2(n23), .A3(opv1[15]), .A4(n102), .Y(n115)
         );
  INVX1_LVT U92 ( .A(opv2[13]), .Y(n99) );
  OR2X1_LVT U93 ( .A1(n99), .A2(opv1[13]), .Y(n22) );
  INVX1_LVT U94 ( .A(opv2[12]), .Y(n29) );
  AO22X1_LVT U95 ( .A1(opv1[12]), .A2(n29), .A3(opv1[13]), .A4(n99), .Y(n110)
         );
  NAND3X0_LVT U96 ( .A1(n115), .A2(n22), .A3(n110), .Y(n33) );
  NOR2X0_LVT U97 ( .A1(n102), .A2(opv1[15]), .Y(n31) );
  AOI22X1_LVT U98 ( .A1(n102), .A2(opv1[15]), .A3(n23), .A4(opv1[14]), .Y(n111) );
  INVX1_LVT U99 ( .A(opv2[11]), .Y(n103) );
  NOR2X0_LVT U100 ( .A1(n103), .A2(opv1[11]), .Y(n28) );
  INVX1_LVT U101 ( .A(opv2[10]), .Y(n24) );
  AOI22X1_LVT U102 ( .A1(n24), .A2(opv1[10]), .A3(n103), .A4(opv1[11]), .Y(
        n106) );
  INVX1_LVT U103 ( .A(opv1[9]), .Y(n25) );
  INVX1_LVT U104 ( .A(opv1[8]), .Y(n34) );
  OA22X1_LVT U105 ( .A1(opv2[9]), .A2(n25), .A3(opv2[8]), .A4(n34), .Y(n27) );
  OA22X1_LVT U106 ( .A1(opv1[11]), .A2(n103), .A3(opv1[10]), .A4(n24), .Y(n109) );
  NAND2X0_LVT U107 ( .A1(opv2[9]), .A2(n25), .Y(n26) );
  NAND2X0_LVT U108 ( .A1(n109), .A2(n26), .Y(n36) );
  OA22X1_LVT U109 ( .A1(n28), .A2(n106), .A3(n27), .A4(n36), .Y(n30) );
  OA22X1_LVT U110 ( .A1(opv1[13]), .A2(n99), .A3(opv1[12]), .A4(n29), .Y(n98)
         );
  NAND2X0_LVT U111 ( .A1(n98), .A2(n115), .Y(n37) );
  OA22X1_LVT U112 ( .A1(n31), .A2(n111), .A3(n30), .A4(n37), .Y(n32) );
  AND2X1_LVT U113 ( .A1(n33), .A2(n32), .Y(n51) );
  AND2X1_LVT U114 ( .A1(opv2[8]), .A2(n34), .Y(n35) );
  OR3X1_LVT U115 ( .A1(n37), .A2(n36), .A3(n35), .Y(n222) );
  INVX1_LVT U116 ( .A(opv2[6]), .Y(n46) );
  INVX1_LVT U117 ( .A(opv2[7]), .Y(n138) );
  OA22X1_LVT U118 ( .A1(opv1[6]), .A2(n46), .A3(opv1[7]), .A4(n138), .Y(n210)
         );
  INVX1_LVT U119 ( .A(opv2[4]), .Y(n43) );
  INVX1_LVT U120 ( .A(opv2[5]), .Y(n134) );
  OA22X1_LVT U121 ( .A1(opv1[4]), .A2(n43), .A3(opv1[5]), .A4(n134), .Y(n219)
         );
  INVX1_LVT U122 ( .A(opv1[1]), .Y(n127) );
  INVX1_LVT U123 ( .A(opv2[3]), .Y(n130) );
  INVX1_LVT U124 ( .A(opv2[2]), .Y(n39) );
  OAI22X1_LVT U125 ( .A1(opv1[3]), .A2(n130), .A3(opv1[2]), .A4(n39), .Y(n131)
         );
  AO21X1_LVT U126 ( .A1(n127), .A2(opv2[1]), .A3(n131), .Y(n199) );
  INVX1_LVT U127 ( .A(n199), .Y(n42) );
  INVX1_LVT U128 ( .A(opv1[0]), .Y(n126) );
  OR2X1_LVT U129 ( .A1(n127), .A2(opv2[1]), .Y(n38) );
  NAND3X0_LVT U130 ( .A1(opv2[0]), .A2(n126), .A3(n38), .Y(n41) );
  OR2X1_LVT U131 ( .A1(n130), .A2(opv1[3]), .Y(n40) );
  AO22X1_LVT U132 ( .A1(opv1[2]), .A2(n39), .A3(opv1[3]), .A4(n130), .Y(n124)
         );
  AO22X1_LVT U133 ( .A1(n42), .A2(n41), .A3(n40), .A4(n124), .Y(n45) );
  OR2X1_LVT U134 ( .A1(n134), .A2(opv1[5]), .Y(n44) );
  AO22X1_LVT U135 ( .A1(opv1[5]), .A2(n134), .A3(opv1[4]), .A4(n43), .Y(n123)
         );
  AO22X1_LVT U136 ( .A1(n219), .A2(n45), .A3(n44), .A4(n123), .Y(n48) );
  OR2X1_LVT U137 ( .A1(n138), .A2(opv1[7]), .Y(n47) );
  AO22X1_LVT U138 ( .A1(opv1[7]), .A2(n138), .A3(opv1[6]), .A4(n46), .Y(n122)
         );
  AOI22X1_LVT U139 ( .A1(n210), .A2(n48), .A3(n47), .A4(n122), .Y(n49) );
  OR2X1_LVT U140 ( .A1(n222), .A2(n49), .Y(n50) );
  AND2X1_LVT U141 ( .A1(n51), .A2(n50), .Y(n62) );
  INVX1_LVT U143 ( .A(opv1[23]), .Y(n147) );
  AO22X1_LVT U144 ( .A1(n831), .A2(opv2[22]), .A3(n147), .A4(opv2[23]), .Y(n63) );
  INVX1_LVT U145 ( .A(opv2[20]), .Y(n65) );
  NOR2X0_LVT U146 ( .A1(n65), .A2(opv1[20]), .Y(n162) );
  INVX1_LVT U147 ( .A(opv2[21]), .Y(n64) );
  NOR2X0_LVT U148 ( .A1(n64), .A2(opv1[21]), .Y(n163) );
  OR3X1_LVT U149 ( .A1(n63), .A2(n162), .A3(n163), .Y(n60) );
  INVX1_LVT U150 ( .A(n60), .Y(n53) );
  INVX1_LVT U151 ( .A(opv2[17]), .Y(n152) );
  INVX1_LVT U152 ( .A(opv1[19]), .Y(n154) );
  INVX1_LVT U153 ( .A(opv1[18]), .Y(n54) );
  AOI22X1_LVT U154 ( .A1(n154), .A2(opv2[19]), .A3(n54), .A4(opv2[18]), .Y(
        n156) );
  OA21X1_LVT U155 ( .A1(opv1[17]), .A2(n152), .A3(n156), .Y(n56) );
  NAND2X0_LVT U157 ( .A1(opv2[16]), .A2(n829), .Y(n52) );
  NAND3X0_LVT U158 ( .A1(n53), .A2(n56), .A3(n52), .Y(n221) );
  AND2X1_LVT U159 ( .A1(opv2[19]), .A2(n154), .Y(n59) );
  OA22X1_LVT U160 ( .A1(opv2[19]), .A2(n154), .A3(opv2[18]), .A4(n54), .Y(n145) );
  OA22X1_LVT U162 ( .A1(opv2[16]), .A2(n829), .A3(opv2[17]), .A4(n830), .Y(n58) );
  INVX1_LVT U163 ( .A(n56), .Y(n57) );
  OA22X1_LVT U164 ( .A1(n59), .A2(n145), .A3(n58), .A4(n57), .Y(n61) );
  OA22X1_LVT U165 ( .A1(n62), .A2(n221), .A3(n61), .A4(n60), .Y(n72) );
  INVX1_LVT U166 ( .A(n63), .Y(n68) );
  INVX1_LVT U167 ( .A(n163), .Y(n67) );
  NAND2X0_LVT U168 ( .A1(opv1[21]), .A2(n64), .Y(n164) );
  NAND2X0_LVT U169 ( .A1(opv1[20]), .A2(n65), .Y(n148) );
  NAND2X0_LVT U170 ( .A1(n164), .A2(n148), .Y(n66) );
  NAND3X0_LVT U171 ( .A1(n68), .A2(n67), .A3(n66), .Y(n71) );
  OR2X1_LVT U172 ( .A1(n147), .A2(opv2[23]), .Y(n169) );
  NAND2X0_LVT U173 ( .A1(opv2[23]), .A2(n147), .Y(n173) );
  INVX1_LVT U174 ( .A(opv2[22]), .Y(n69) );
  NAND3X0_LVT U175 ( .A1(opv1[22]), .A2(n173), .A3(n69), .Y(n70) );
  AND4X1_LVT U176 ( .A1(n72), .A2(n71), .A3(n169), .A4(n70), .Y(n75) );
  AND2X1_LVT U177 ( .A1(opv2[27]), .A2(n175), .Y(n74) );
  OA22X1_LVT U178 ( .A1(opv2[26]), .A2(n73), .A3(opv2[27]), .A4(n175), .Y(n93)
         );
  OA222X1_LVT U179 ( .A1(n77), .A2(n76), .A3(n198), .A4(n75), .A5(n74), .A6(
        n93), .Y(n83) );
  NAND2X0_LVT U180 ( .A1(opv2[28]), .A2(n78), .Y(n91) );
  NAND2X0_LVT U181 ( .A1(opv2[29]), .A2(n79), .Y(n80) );
  NAND2X0_LVT U182 ( .A1(n91), .A2(n80), .Y(n200) );
  INVX1_LVT U183 ( .A(opv2[31]), .Y(n82) );
  OR2X1_LVT U184 ( .A1(n82), .A2(opv1[31]), .Y(n202) );
  INVX1_LVT U185 ( .A(opv2[30]), .Y(n87) );
  OR2X1_LVT U186 ( .A1(n87), .A2(opv1[30]), .Y(n201) );
  NAND2X0_LVT U187 ( .A1(n202), .A2(n201), .Y(n81) );
  AO221X1_LVT U188 ( .A1(n85), .A2(n83), .A3(n85), .A4(n200), .A5(n81), .Y(n90) );
  NAND2X0_LVT U189 ( .A1(opv1[31]), .A2(n82), .Y(n206) );
  NAND2X0_LVT U190 ( .A1(n201), .A2(n206), .Y(n86) );
  OR2X1_LVT U191 ( .A1(n200), .A2(n83), .Y(n84) );
  OA221X1_LVT U192 ( .A1(n86), .A2(n85), .A3(n86), .A4(n84), .A5(n202), .Y(n88) );
  NAND2X0_LVT U193 ( .A1(n202), .A2(n206), .Y(n190) );
  NAND2X0_LVT U194 ( .A1(opv1[30]), .A2(n87), .Y(n205) );
  OA22X1_LVT U195 ( .A1(inst[13]), .A2(n88), .A3(n190), .A4(n205), .Y(n89) );
  OA221X1_LVT U196 ( .A1(n836), .A2(n90), .A3(n836), .A4(n206), .A5(n89), .Y(
        n195) );
  INVX1_LVT U197 ( .A(opv2[29]), .Y(n181) );
  AO222X1_LVT U198 ( .A1(opv1[29]), .A2(n91), .A3(opv1[29]), .A4(n181), .A5(
        n91), .A6(n181), .Y(n187) );
  INVX1_LVT U199 ( .A(opv2[25]), .Y(n94) );
  NAND2X0_LVT U200 ( .A1(opv1[25]), .A2(n94), .Y(n92) );
  NAND2X0_LVT U201 ( .A1(n93), .A2(n92), .Y(n180) );
  INVX1_LVT U202 ( .A(opv2[24]), .Y(n95) );
  OA22X1_LVT U203 ( .A1(opv1[24]), .A2(n95), .A3(opv1[25]), .A4(n94), .Y(n179)
         );
  INVX1_LVT U204 ( .A(n180), .Y(n97) );
  NAND2X0_LVT U205 ( .A1(opv1[24]), .A2(n95), .Y(n96) );
  NAND2X0_LVT U206 ( .A1(n97), .A2(n96), .Y(n197) );
  INVX1_LVT U207 ( .A(n98), .Y(n101) );
  NAND2X0_LVT U208 ( .A1(opv1[13]), .A2(n99), .Y(n100) );
  NAND3X0_LVT U209 ( .A1(n111), .A2(n101), .A3(n100), .Y(n117) );
  AND2X1_LVT U210 ( .A1(opv1[15]), .A2(n102), .Y(n114) );
  AND2X1_LVT U211 ( .A1(opv1[11]), .A2(n103), .Y(n108) );
  INVX1_LVT U212 ( .A(opv2[8]), .Y(n118) );
  INVX1_LVT U213 ( .A(opv2[9]), .Y(n104) );
  OA22X1_LVT U214 ( .A1(opv1[8]), .A2(n118), .A3(opv1[9]), .A4(n104), .Y(n107)
         );
  NAND2X0_LVT U215 ( .A1(opv1[9]), .A2(n104), .Y(n105) );
  NAND2X0_LVT U216 ( .A1(n106), .A2(n105), .Y(n120) );
  OA22X1_LVT U217 ( .A1(n109), .A2(n108), .A3(n107), .A4(n120), .Y(n113) );
  INVX1_LVT U218 ( .A(n110), .Y(n112) );
  NAND2X0_LVT U219 ( .A1(n112), .A2(n111), .Y(n121) );
  OA22X1_LVT U220 ( .A1(n115), .A2(n114), .A3(n113), .A4(n121), .Y(n116) );
  AND2X1_LVT U221 ( .A1(n117), .A2(n116), .Y(n144) );
  AND2X1_LVT U222 ( .A1(opv1[8]), .A2(n118), .Y(n119) );
  OR3X1_LVT U223 ( .A1(n121), .A2(n120), .A3(n119), .Y(n214) );
  INVX1_LVT U224 ( .A(n122), .Y(n211) );
  INVX1_LVT U225 ( .A(n123), .Y(n218) );
  INVX1_LVT U226 ( .A(n124), .Y(n125) );
  OA21X1_LVT U227 ( .A1(opv2[1]), .A2(n127), .A3(n125), .Y(n209) );
  NAND2X0_LVT U228 ( .A1(opv2[0]), .A2(n126), .Y(n129) );
  NAND2X0_LVT U229 ( .A1(opv2[1]), .A2(n127), .Y(n128) );
  NAND2X0_LVT U230 ( .A1(n129), .A2(n128), .Y(n133) );
  NAND2X0_LVT U231 ( .A1(opv1[3]), .A2(n130), .Y(n132) );
  AO22X1_LVT U232 ( .A1(n209), .A2(n133), .A3(n132), .A4(n131), .Y(n137) );
  INVX1_LVT U233 ( .A(n219), .Y(n136) );
  NAND2X0_LVT U234 ( .A1(opv1[5]), .A2(n134), .Y(n135) );
  AO22X1_LVT U235 ( .A1(n218), .A2(n137), .A3(n136), .A4(n135), .Y(n141) );
  NAND2X0_LVT U236 ( .A1(opv1[7]), .A2(n138), .Y(n140) );
  INVX1_LVT U237 ( .A(n210), .Y(n139) );
  AOI22X1_LVT U238 ( .A1(n211), .A2(n141), .A3(n140), .A4(n139), .Y(n142) );
  OR2X1_LVT U239 ( .A1(n214), .A2(n142), .Y(n143) );
  AND2X1_LVT U240 ( .A1(n144), .A2(n143), .Y(n161) );
  OA21X1_LVT U241 ( .A1(opv2[17]), .A2(n830), .A3(n145), .Y(n153) );
  OA22X1_LVT U242 ( .A1(opv2[23]), .A2(n147), .A3(opv2[22]), .A4(n831), .Y(
        n165) );
  NAND3X0_LVT U243 ( .A1(n165), .A2(n164), .A3(n148), .Y(n159) );
  INVX1_LVT U244 ( .A(n159), .Y(n150) );
  INVX1_LVT U245 ( .A(opv2[16]), .Y(n151) );
  NAND2X0_LVT U246 ( .A1(opv1[16]), .A2(n151), .Y(n149) );
  NAND3X0_LVT U247 ( .A1(n153), .A2(n150), .A3(n149), .Y(n213) );
  OA22X1_LVT U248 ( .A1(opv1[17]), .A2(n152), .A3(opv1[16]), .A4(n151), .Y(
        n158) );
  INVX1_LVT U249 ( .A(n153), .Y(n157) );
  NOR2X0_LVT U250 ( .A1(n154), .A2(opv2[19]), .Y(n155) );
  OA22X1_LVT U251 ( .A1(n158), .A2(n157), .A3(n156), .A4(n155), .Y(n160) );
  OA22X1_LVT U252 ( .A1(n161), .A2(n213), .A3(n160), .A4(n159), .Y(n174) );
  INVX1_LVT U253 ( .A(n162), .Y(n168) );
  INVX1_LVT U254 ( .A(n163), .Y(n167) );
  NAND2X0_LVT U255 ( .A1(n165), .A2(n164), .Y(n166) );
  AO21X1_LVT U256 ( .A1(n168), .A2(n167), .A3(n166), .Y(n172) );
  NAND3X0_LVT U257 ( .A1(opv2[22]), .A2(n831), .A3(n169), .Y(n171) );
  AND4X1_LVT U258 ( .A1(n174), .A2(n173), .A3(n172), .A4(n171), .Y(n178) );
  NOR2X0_LVT U259 ( .A1(n175), .A2(opv2[27]), .Y(n176) );
  OA222X1_LVT U260 ( .A1(n180), .A2(n179), .A3(n197), .A4(n178), .A5(n177), 
        .A6(n176), .Y(n186) );
  NAND2X0_LVT U261 ( .A1(opv1[29]), .A2(n181), .Y(n183) );
  NAND2X0_LVT U262 ( .A1(n183), .A2(n182), .Y(n204) );
  NAND2X0_LVT U263 ( .A1(n206), .A2(n205), .Y(n184) );
  AO221X1_LVT U264 ( .A1(n187), .A2(n186), .A3(n187), .A4(n204), .A5(n184), 
        .Y(n193) );
  INVX1_LVT U265 ( .A(n202), .Y(n189) );
  INVX1_LVT U266 ( .A(n205), .Y(n185) );
  AO221X1_LVT U267 ( .A1(n187), .A2(n186), .A3(n187), .A4(n204), .A5(n185), 
        .Y(n188) );
  OA21X1_LVT U268 ( .A1(n189), .A2(n188), .A3(n206), .Y(n191) );
  OA22X1_LVT U269 ( .A1(inst[13]), .A2(n191), .A3(n190), .A4(n201), .Y(n192)
         );
  OA221X1_LVT U270 ( .A1(n836), .A2(n193), .A3(n836), .A4(n202), .A5(n192), 
        .Y(n194) );
  AO221X1_LVT U271 ( .A1(inst[12]), .A2(n195), .A3(n813), .A4(n194), .A5(n812), 
        .Y(n225) );
  NAND2X0_LVT U272 ( .A1(n812), .A2(n836), .Y(n774) );
  HADDX1_LVT U273 ( .A0(opv1[0]), .B0(opv2[0]), .SO(n196) );
  NOR4X1_LVT U274 ( .A1(n199), .A2(n198), .A3(n197), .A4(n196), .Y(n217) );
  INVX1_LVT U275 ( .A(n200), .Y(n203) );
  NAND3X0_LVT U276 ( .A1(n203), .A2(n202), .A3(n201), .Y(n215) );
  INVX1_LVT U277 ( .A(n204), .Y(n207) );
  AND3X1_LVT U278 ( .A1(n207), .A2(n206), .A3(n205), .Y(n208) );
  NAND4X0_LVT U279 ( .A1(n211), .A2(n210), .A3(n209), .A4(n208), .Y(n212) );
  NOR4X1_LVT U280 ( .A1(n215), .A2(n214), .A3(n213), .A4(n212), .Y(n216) );
  NAND4X0_LVT U281 ( .A1(n219), .A2(n218), .A3(n217), .A4(n216), .Y(n220) );
  OR3X1_LVT U282 ( .A1(n222), .A2(n221), .A3(n220), .Y(n223) );
  HADDX1_LVT U283 ( .A0(inst[12]), .B0(n223), .SO(n224) );
  AO221X1_LVT U284 ( .A1(n225), .A2(n774), .A3(n225), .A4(n224), .A5(n780), 
        .Y(n226) );
  NAND2X0_LVT U286 ( .A1(inst[15]), .A2(n227), .Y(n589) );
  INVX1_LVT U287 ( .A(n589), .Y(reg_addr1[0]) );
  INVX1_LVT U288 ( .A(ex_aluop[3]), .Y(n228) );
  NOR3X0_LVT U289 ( .A1(ex_aluop[0]), .A2(ex_aluop[1]), .A3(n228), .Y(n230) );
  OA221X1_LVT U291 ( .A1(ex_aluop[2]), .A2(n230), .A3(n810), .A4(n228), .A5(
        ex_aluop[4]), .Y(n253) );
  HADDX1_LVT U292 ( .A0(ex_reg_waddr[0]), .B0(reg_addr1[0]), .SO(n236) );
  INVX1_LVT U293 ( .A(re1), .Y(n235) );
  OAI22X1_LVT U294 ( .A1(n581), .A2(ex_reg_waddr[4]), .A3(n588), .A4(
        ex_reg_waddr[3]), .Y(n231) );
  AO221X1_LVT U295 ( .A1(n581), .A2(ex_reg_waddr[4]), .A3(n588), .A4(
        ex_reg_waddr[3]), .A5(n231), .Y(n234) );
  OAI22X1_LVT U296 ( .A1(n582), .A2(ex_reg_waddr[2]), .A3(n583), .A4(
        ex_reg_waddr[1]), .Y(n232) );
  AO221X1_LVT U297 ( .A1(n582), .A2(ex_reg_waddr[2]), .A3(n583), .A4(
        ex_reg_waddr[1]), .A5(n232), .Y(n233) );
  NOR4X1_LVT U298 ( .A1(n236), .A2(n235), .A3(n234), .A4(n233), .Y(n579) );
  AND2X1_LVT U302 ( .A1(inst[21]), .A2(n243), .Y(reg_addr2[1]) );
  AND3X1_LVT U303 ( .A1(n492), .A2(n238), .A3(n269), .Y(n241) );
  AO21X1_LVT U304 ( .A1(n241), .A2(n240), .A3(n239), .Y(n242) );
  NAND2X0_LVT U305 ( .A1(n751), .A2(n242), .Y(n752) );
  AND2X2_LVT U308 ( .A1(inst[24]), .A2(n243), .Y(reg_addr2[4]) );
  HADDX1_LVT U309 ( .A0(ex_reg_waddr[4]), .B0(reg_addr2[4]), .SO(n251) );
  OAI22X1_LVT U311 ( .A1(n246), .A2(ex_reg_waddr[3]), .A3(n815), .A4(
        ex_reg_waddr[1]), .Y(n244) );
  AO221X1_LVT U312 ( .A1(n246), .A2(ex_reg_waddr[3]), .A3(n815), .A4(
        ex_reg_waddr[1]), .A5(n244), .Y(n250) );
  OAI22X1_LVT U313 ( .A1(n248), .A2(ex_reg_waddr[0]), .A3(n260), .A4(
        ex_reg_waddr[2]), .Y(n247) );
  AO221X1_LVT U314 ( .A1(n248), .A2(ex_reg_waddr[0]), .A3(n260), .A4(
        ex_reg_waddr[2]), .A5(n247), .Y(n249) );
  NOR4X1_LVT U315 ( .A1(n252), .A2(n251), .A3(n250), .A4(n249), .Y(n258) );
  NAND2X0_LVT U319 ( .A1(n237), .A2(n254), .Y(stallreq) );
  NAND2X0_LVT U327 ( .A1(ex_we), .A2(n258), .Y(n272) );
  INVX1_LVT U328 ( .A(mem_reg_waddr[0]), .Y(n586) );
  AOI22X1_LVT U329 ( .A1(n586), .A2(reg_addr2[0]), .A3(n260), .A4(
        mem_reg_waddr[2]), .Y(n259) );
  OA221X1_LVT U330 ( .A1(n586), .A2(reg_addr2[0]), .A3(n260), .A4(
        mem_reg_waddr[2]), .A5(n259), .Y(n266) );
  INVX1_LVT U332 ( .A(mem_reg_waddr[4]), .Y(n261) );
  OA221X1_LVT U333 ( .A1(mem_reg_waddr[4]), .A2(n818), .A3(n261), .A4(inst[24]), .A5(re2), .Y(n265) );
  INVX1_LVT U334 ( .A(mem_reg_waddr[3]), .Y(n585) );
  INVX1_LVT U335 ( .A(mem_reg_waddr[1]), .Y(n584) );
  AOI22X1_LVT U336 ( .A1(n585), .A2(reg_addr2[3]), .A3(n584), .A4(reg_addr2[1]), .Y(n263) );
  OA221X1_LVT U337 ( .A1(n585), .A2(reg_addr2[3]), .A3(n584), .A4(reg_addr2[1]), .A5(n263), .Y(n264) );
  NAND4X0_LVT U338 ( .A1(mem_we), .A2(n266), .A3(n265), .A4(n264), .Y(n271) );
  AO22X1_LVT U342 ( .A1(ex_reg_wdata[11]), .A2(n257), .A3(n267), .A4(
        reg_data2[11]), .Y(n268) );
  INVX1_LVT U343 ( .A(n268), .Y(n277) );
  NAND3X0_LVT U344 ( .A1(n751), .A2(inst[2]), .A3(n748), .Y(n739) );
  NAND2X0_LVT U348 ( .A1(inst[12]), .A2(n836), .Y(n759) );
  AND3X2_LVT U349 ( .A1(n765), .A2(n269), .A3(n759), .Y(n749) );
  AO22X1_LVT U350 ( .A1(pc[11]), .A2(n665), .A3(inst[31]), .A4(n749), .Y(n270)
         );
  INVX1_LVT U351 ( .A(n270), .Y(n276) );
  INVX1_LVT U352 ( .A(n271), .Y(n273) );
  NAND2X0_LVT U356 ( .A1(mem_reg_wdata[11]), .A2(n274), .Y(n275) );
  NAND3X0_LVT U357 ( .A1(n277), .A2(n276), .A3(n275), .Y(N707) );
  AO22X1_LVT U358 ( .A1(ex_reg_wdata[10]), .A2(n257), .A3(mem_reg_wdata[10]), 
        .A4(n274), .Y(n278) );
  INVX1_LVT U359 ( .A(n278), .Y(n282) );
  AO22X1_LVT U360 ( .A1(n834), .A2(n665), .A3(inst[30]), .A4(n749), .Y(n279)
         );
  INVX1_LVT U361 ( .A(n279), .Y(n281) );
  NAND2X0_LVT U362 ( .A1(n267), .A2(reg_data2[10]), .Y(n280) );
  NAND3X0_LVT U363 ( .A1(n282), .A2(n281), .A3(n280), .Y(N706) );
  AO22X1_LVT U364 ( .A1(ex_reg_wdata[9]), .A2(n257), .A3(mem_reg_wdata[9]), 
        .A4(n274), .Y(n283) );
  INVX1_LVT U365 ( .A(n283), .Y(n287) );
  AO22X1_LVT U366 ( .A1(pc[9]), .A2(n665), .A3(inst[29]), .A4(n749), .Y(n284)
         );
  INVX1_LVT U367 ( .A(n284), .Y(n286) );
  NAND2X0_LVT U368 ( .A1(n267), .A2(reg_data2[9]), .Y(n285) );
  NAND3X0_LVT U369 ( .A1(n287), .A2(n286), .A3(n285), .Y(N705) );
  AO22X1_LVT U370 ( .A1(ex_reg_wdata[8]), .A2(n257), .A3(mem_reg_wdata[8]), 
        .A4(n274), .Y(n288) );
  INVX1_LVT U371 ( .A(n288), .Y(n292) );
  AO22X1_LVT U372 ( .A1(pc[8]), .A2(n665), .A3(inst[28]), .A4(n749), .Y(n289)
         );
  INVX1_LVT U373 ( .A(n289), .Y(n291) );
  NAND2X0_LVT U374 ( .A1(n267), .A2(reg_data2[8]), .Y(n290) );
  NAND3X0_LVT U375 ( .A1(n292), .A2(n291), .A3(n290), .Y(N704) );
  AO22X1_LVT U376 ( .A1(ex_reg_wdata[7]), .A2(n257), .A3(mem_reg_wdata[7]), 
        .A4(n274), .Y(n293) );
  INVX1_LVT U377 ( .A(n293), .Y(n297) );
  AO22X1_LVT U378 ( .A1(pc[7]), .A2(n665), .A3(inst[27]), .A4(n749), .Y(n294)
         );
  INVX1_LVT U379 ( .A(n294), .Y(n296) );
  NAND2X0_LVT U380 ( .A1(n267), .A2(reg_data2[7]), .Y(n295) );
  NAND3X0_LVT U381 ( .A1(n297), .A2(n296), .A3(n295), .Y(N703) );
  AO22X1_LVT U382 ( .A1(ex_reg_wdata[6]), .A2(n257), .A3(mem_reg_wdata[6]), 
        .A4(n274), .Y(n298) );
  INVX1_LVT U383 ( .A(n298), .Y(n302) );
  AO22X1_LVT U384 ( .A1(pc[6]), .A2(n665), .A3(inst[26]), .A4(n749), .Y(n299)
         );
  INVX1_LVT U385 ( .A(n299), .Y(n301) );
  NAND2X0_LVT U386 ( .A1(n267), .A2(reg_data2[6]), .Y(n300) );
  NAND3X0_LVT U387 ( .A1(n302), .A2(n301), .A3(n300), .Y(N702) );
  AO22X1_LVT U388 ( .A1(ex_reg_wdata[5]), .A2(n257), .A3(mem_reg_wdata[5]), 
        .A4(n274), .Y(n303) );
  INVX1_LVT U389 ( .A(n303), .Y(n307) );
  AO22X1_LVT U390 ( .A1(pc[5]), .A2(n665), .A3(inst[25]), .A4(n749), .Y(n304)
         );
  INVX1_LVT U391 ( .A(n304), .Y(n306) );
  NAND2X0_LVT U392 ( .A1(n267), .A2(reg_data2[5]), .Y(n305) );
  NAND3X0_LVT U393 ( .A1(n307), .A2(n306), .A3(n305), .Y(N701) );
  AO22X1_LVT U394 ( .A1(ex_reg_wdata[4]), .A2(n257), .A3(n267), .A4(
        reg_data2[4]), .Y(n308) );
  INVX1_LVT U395 ( .A(n308), .Y(n313) );
  INVX1_LVT U396 ( .A(n309), .Y(n331) );
  AO22X1_LVT U397 ( .A1(pc[4]), .A2(n665), .A3(n331), .A4(inst[24]), .Y(n310)
         );
  INVX1_LVT U398 ( .A(n310), .Y(n312) );
  NAND2X0_LVT U399 ( .A1(mem_reg_wdata[4]), .A2(n274), .Y(n311) );
  NAND3X0_LVT U400 ( .A1(n313), .A2(n312), .A3(n311), .Y(N700) );
  AO22X1_LVT U401 ( .A1(ex_reg_wdata[3]), .A2(n257), .A3(n267), .A4(
        reg_data2[3]), .Y(n314) );
  INVX1_LVT U402 ( .A(n314), .Y(n318) );
  AO22X1_LVT U403 ( .A1(pc[3]), .A2(n665), .A3(n331), .A4(inst[23]), .Y(n315)
         );
  INVX1_LVT U404 ( .A(n315), .Y(n317) );
  NAND2X0_LVT U405 ( .A1(mem_reg_wdata[3]), .A2(n274), .Y(n316) );
  NAND3X0_LVT U406 ( .A1(n318), .A2(n317), .A3(n316), .Y(N699) );
  AO22X1_LVT U407 ( .A1(ex_reg_wdata[2]), .A2(n257), .A3(n267), .A4(
        reg_data2[2]), .Y(n319) );
  INVX1_LVT U408 ( .A(n319), .Y(n323) );
  AO22X1_LVT U409 ( .A1(pc[2]), .A2(n665), .A3(n331), .A4(inst[22]), .Y(n320)
         );
  INVX1_LVT U410 ( .A(n320), .Y(n322) );
  NAND2X0_LVT U411 ( .A1(mem_reg_wdata[2]), .A2(n274), .Y(n321) );
  NAND3X0_LVT U412 ( .A1(n323), .A2(n322), .A3(n321), .Y(N698) );
  AO22X1_LVT U414 ( .A1(ex_reg_wdata[1]), .A2(n257), .A3(n267), .A4(
        reg_data2[1]), .Y(n324) );
  INVX1_LVT U415 ( .A(n324), .Y(n328) );
  AO22X1_LVT U416 ( .A1(n331), .A2(inst[21]), .A3(n665), .A4(pc[1]), .Y(n325)
         );
  INVX1_LVT U417 ( .A(n325), .Y(n327) );
  NAND2X0_LVT U418 ( .A1(mem_reg_wdata[1]), .A2(n274), .Y(n326) );
  NAND3X0_LVT U419 ( .A1(n328), .A2(n327), .A3(n326), .Y(N697) );
  AO22X1_LVT U420 ( .A1(ex_reg_wdata[0]), .A2(n257), .A3(n267), .A4(
        reg_data2[0]), .Y(n330) );
  INVX1_LVT U421 ( .A(n330), .Y(n335) );
  AO22X1_LVT U422 ( .A1(n331), .A2(inst[20]), .A3(pc[0]), .A4(n665), .Y(n332)
         );
  INVX1_LVT U423 ( .A(n332), .Y(n334) );
  NAND2X0_LVT U424 ( .A1(mem_reg_wdata[0]), .A2(n274), .Y(n333) );
  NAND3X0_LVT U425 ( .A1(n335), .A2(n334), .A3(n333), .Y(N696) );
  NAND4X0_LVT U426 ( .A1(pc[2]), .A2(pc[3]), .A3(pc[4]), .A4(pc[5]), .Y(n436)
         );
  INVX1_LVT U427 ( .A(n436), .Y(n433) );
  NAND2X0_LVT U428 ( .A1(n433), .A2(pc[6]), .Y(n432) );
  INVX1_LVT U429 ( .A(n432), .Y(n429) );
  NAND2X0_LVT U430 ( .A1(n429), .A2(pc[7]), .Y(n428) );
  INVX1_LVT U431 ( .A(n428), .Y(n425) );
  NAND2X0_LVT U432 ( .A1(n425), .A2(pc[8]), .Y(n424) );
  INVX1_LVT U433 ( .A(n424), .Y(n421) );
  NAND2X0_LVT U434 ( .A1(n421), .A2(pc[9]), .Y(n420) );
  INVX1_LVT U435 ( .A(n420), .Y(n417) );
  NAND2X0_LVT U436 ( .A1(n417), .A2(pc[10]), .Y(n416) );
  INVX1_LVT U437 ( .A(n416), .Y(n413) );
  NAND2X0_LVT U438 ( .A1(n413), .A2(pc[11]), .Y(n412) );
  INVX1_LVT U439 ( .A(n412), .Y(n409) );
  NAND2X0_LVT U440 ( .A1(n409), .A2(pc[12]), .Y(n408) );
  INVX1_LVT U441 ( .A(n408), .Y(n405) );
  NAND2X0_LVT U442 ( .A1(n405), .A2(pc[13]), .Y(n404) );
  INVX1_LVT U443 ( .A(n404), .Y(n401) );
  NAND2X0_LVT U444 ( .A1(n401), .A2(pc[14]), .Y(n400) );
  INVX1_LVT U445 ( .A(n400), .Y(n397) );
  NAND2X0_LVT U446 ( .A1(n397), .A2(pc[15]), .Y(n396) );
  INVX1_LVT U447 ( .A(n396), .Y(n393) );
  NAND2X0_LVT U448 ( .A1(n393), .A2(pc[16]), .Y(n392) );
  INVX1_LVT U449 ( .A(n392), .Y(n389) );
  NAND2X0_LVT U450 ( .A1(n389), .A2(pc[17]), .Y(n388) );
  INVX1_LVT U451 ( .A(n388), .Y(n385) );
  NAND2X0_LVT U452 ( .A1(n385), .A2(pc[18]), .Y(n384) );
  INVX1_LVT U453 ( .A(n384), .Y(n381) );
  NAND2X0_LVT U454 ( .A1(n381), .A2(pc[19]), .Y(n380) );
  INVX1_LVT U455 ( .A(n380), .Y(n377) );
  NAND2X0_LVT U456 ( .A1(n377), .A2(pc[20]), .Y(n376) );
  INVX1_LVT U457 ( .A(n376), .Y(n373) );
  NAND2X0_LVT U458 ( .A1(n373), .A2(pc[21]), .Y(n372) );
  INVX1_LVT U459 ( .A(n372), .Y(n369) );
  NAND2X0_LVT U460 ( .A1(n369), .A2(pc[22]), .Y(n368) );
  INVX1_LVT U461 ( .A(n368), .Y(n365) );
  NAND2X0_LVT U462 ( .A1(n365), .A2(pc[23]), .Y(n364) );
  INVX1_LVT U463 ( .A(n364), .Y(n360) );
  NAND2X0_LVT U464 ( .A1(n360), .A2(pc[24]), .Y(n359) );
  INVX1_LVT U465 ( .A(n359), .Y(n356) );
  NAND2X0_LVT U466 ( .A1(n356), .A2(pc[25]), .Y(n355) );
  INVX1_LVT U467 ( .A(n355), .Y(n352) );
  NAND2X0_LVT U468 ( .A1(n352), .A2(pc[26]), .Y(n351) );
  INVX1_LVT U469 ( .A(n351), .Y(n348) );
  NAND2X0_LVT U470 ( .A1(n348), .A2(pc[27]), .Y(n347) );
  INVX1_LVT U471 ( .A(n347), .Y(n344) );
  NAND2X0_LVT U472 ( .A1(n344), .A2(pc[28]), .Y(n343) );
  INVX1_LVT U473 ( .A(n343), .Y(n340) );
  NAND2X0_LVT U474 ( .A1(n340), .A2(pc[29]), .Y(n339) );
  INVX1_LVT U475 ( .A(n339), .Y(n336) );
  NAND2X0_LVT U476 ( .A1(n336), .A2(pc[30]), .Y(n728) );
  AND2X1_LVT U479 ( .A1(n728), .A2(n821), .Y(n338) );
  OR2X1_LVT U480 ( .A1(pc[30]), .A2(n336), .Y(n337) );
  AND2X1_LVT U481 ( .A1(n338), .A2(n337), .Y(link_addr[30]) );
  AND2X1_LVT U482 ( .A1(n339), .A2(n821), .Y(n342) );
  OR2X1_LVT U483 ( .A1(pc[29]), .A2(n340), .Y(n341) );
  AND2X1_LVT U484 ( .A1(n342), .A2(n341), .Y(link_addr[29]) );
  AND2X1_LVT U485 ( .A1(n343), .A2(n821), .Y(n346) );
  OR2X1_LVT U486 ( .A1(pc[28]), .A2(n344), .Y(n345) );
  AND2X1_LVT U487 ( .A1(n346), .A2(n345), .Y(link_addr[28]) );
  AND2X1_LVT U488 ( .A1(n347), .A2(n821), .Y(n350) );
  OR2X1_LVT U489 ( .A1(pc[27]), .A2(n348), .Y(n349) );
  AND2X1_LVT U490 ( .A1(n350), .A2(n349), .Y(link_addr[27]) );
  AND2X1_LVT U491 ( .A1(n351), .A2(n821), .Y(n354) );
  OR2X1_LVT U492 ( .A1(pc[26]), .A2(n352), .Y(n353) );
  AND2X1_LVT U493 ( .A1(n354), .A2(n353), .Y(link_addr[26]) );
  AND2X1_LVT U494 ( .A1(n355), .A2(n821), .Y(n358) );
  OR2X1_LVT U495 ( .A1(pc[25]), .A2(n356), .Y(n357) );
  AND2X1_LVT U496 ( .A1(n358), .A2(n357), .Y(link_addr[25]) );
  AND2X1_LVT U497 ( .A1(n359), .A2(n821), .Y(n362) );
  OR2X1_LVT U498 ( .A1(pc[24]), .A2(n360), .Y(n361) );
  AND2X1_LVT U499 ( .A1(n362), .A2(n361), .Y(link_addr[24]) );
  AND2X1_LVT U501 ( .A1(n364), .A2(n821), .Y(n367) );
  OR2X1_LVT U502 ( .A1(pc[23]), .A2(n365), .Y(n366) );
  AND2X1_LVT U503 ( .A1(n367), .A2(n366), .Y(link_addr[23]) );
  AND2X1_LVT U504 ( .A1(n368), .A2(n821), .Y(n371) );
  OR2X1_LVT U505 ( .A1(pc[22]), .A2(n369), .Y(n370) );
  AND2X1_LVT U506 ( .A1(n371), .A2(n370), .Y(link_addr[22]) );
  AND2X1_LVT U507 ( .A1(n372), .A2(n821), .Y(n375) );
  OR2X1_LVT U508 ( .A1(pc[21]), .A2(n373), .Y(n374) );
  AND2X1_LVT U509 ( .A1(n375), .A2(n374), .Y(link_addr[21]) );
  AND2X1_LVT U510 ( .A1(n376), .A2(n821), .Y(n379) );
  OR2X1_LVT U511 ( .A1(pc[20]), .A2(n377), .Y(n378) );
  AND2X1_LVT U512 ( .A1(n379), .A2(n378), .Y(link_addr[20]) );
  AND2X1_LVT U513 ( .A1(n380), .A2(n821), .Y(n383) );
  OR2X1_LVT U514 ( .A1(pc[19]), .A2(n381), .Y(n382) );
  AND2X1_LVT U515 ( .A1(n383), .A2(n382), .Y(link_addr[19]) );
  AND2X1_LVT U516 ( .A1(n384), .A2(n821), .Y(n387) );
  OR2X1_LVT U517 ( .A1(pc[18]), .A2(n385), .Y(n386) );
  AND2X1_LVT U518 ( .A1(n387), .A2(n386), .Y(link_addr[18]) );
  AND2X1_LVT U519 ( .A1(n388), .A2(n821), .Y(n391) );
  OR2X1_LVT U520 ( .A1(pc[17]), .A2(n389), .Y(n390) );
  AND2X1_LVT U521 ( .A1(n391), .A2(n390), .Y(link_addr[17]) );
  AND2X1_LVT U522 ( .A1(n392), .A2(n821), .Y(n395) );
  OR2X1_LVT U523 ( .A1(pc[16]), .A2(n393), .Y(n394) );
  AND2X1_LVT U524 ( .A1(n395), .A2(n394), .Y(link_addr[16]) );
  AND2X1_LVT U525 ( .A1(n396), .A2(n821), .Y(n399) );
  OR2X1_LVT U526 ( .A1(pc[15]), .A2(n397), .Y(n398) );
  AND2X1_LVT U527 ( .A1(n399), .A2(n398), .Y(link_addr[15]) );
  AND2X1_LVT U528 ( .A1(n400), .A2(n821), .Y(n403) );
  OR2X1_LVT U529 ( .A1(pc[14]), .A2(n401), .Y(n402) );
  AND2X1_LVT U530 ( .A1(n403), .A2(n402), .Y(link_addr[14]) );
  AND2X1_LVT U531 ( .A1(n404), .A2(n821), .Y(n407) );
  OR2X1_LVT U532 ( .A1(pc[13]), .A2(n405), .Y(n406) );
  AND2X1_LVT U533 ( .A1(n407), .A2(n406), .Y(link_addr[13]) );
  AND2X1_LVT U534 ( .A1(n408), .A2(n821), .Y(n411) );
  OR2X1_LVT U535 ( .A1(pc[12]), .A2(n409), .Y(n410) );
  AND2X1_LVT U536 ( .A1(n411), .A2(n410), .Y(link_addr[12]) );
  AND2X1_LVT U537 ( .A1(n412), .A2(n821), .Y(n415) );
  OR2X1_LVT U538 ( .A1(pc[11]), .A2(n413), .Y(n414) );
  AND2X1_LVT U539 ( .A1(n415), .A2(n414), .Y(link_addr[11]) );
  AND2X1_LVT U540 ( .A1(n416), .A2(n821), .Y(n419) );
  OR2X1_LVT U541 ( .A1(pc[10]), .A2(n417), .Y(n418) );
  AND2X1_LVT U542 ( .A1(n419), .A2(n418), .Y(link_addr[10]) );
  AND2X1_LVT U543 ( .A1(n420), .A2(n821), .Y(n423) );
  OR2X1_LVT U544 ( .A1(pc[9]), .A2(n421), .Y(n422) );
  AND2X1_LVT U545 ( .A1(n423), .A2(n422), .Y(link_addr[9]) );
  AND2X1_LVT U546 ( .A1(n424), .A2(n821), .Y(n427) );
  OR2X1_LVT U547 ( .A1(pc[8]), .A2(n425), .Y(n426) );
  AND2X1_LVT U548 ( .A1(n427), .A2(n426), .Y(link_addr[8]) );
  AND2X1_LVT U549 ( .A1(n428), .A2(n821), .Y(n431) );
  OR2X1_LVT U550 ( .A1(pc[7]), .A2(n429), .Y(n430) );
  AND2X1_LVT U551 ( .A1(n431), .A2(n430), .Y(link_addr[7]) );
  AND2X1_LVT U552 ( .A1(n432), .A2(n821), .Y(n435) );
  OR2X1_LVT U553 ( .A1(pc[6]), .A2(n433), .Y(n434) );
  AND2X1_LVT U554 ( .A1(n435), .A2(n434), .Y(link_addr[6]) );
  AND2X1_LVT U555 ( .A1(n436), .A2(n821), .Y(n439) );
  NAND3X0_LVT U556 ( .A1(pc[2]), .A2(pc[3]), .A3(pc[4]), .Y(n440) );
  INVX1_LVT U557 ( .A(n440), .Y(n437) );
  OR2X1_LVT U558 ( .A1(pc[5]), .A2(n437), .Y(n438) );
  AND2X1_LVT U559 ( .A1(n439), .A2(n438), .Y(link_addr[5]) );
  AND2X1_LVT U560 ( .A1(n440), .A2(n821), .Y(n443) );
  AND2X1_LVT U561 ( .A1(pc[2]), .A2(pc[3]), .Y(n441) );
  OR2X1_LVT U562 ( .A1(pc[4]), .A2(n441), .Y(n442) );
  AND2X1_LVT U563 ( .A1(n443), .A2(n442), .Y(link_addr[4]) );
  INVX1_LVT U564 ( .A(n492), .Y(n445) );
  AO22X1_LVT U569 ( .A1(n823), .A2(reg_data1[0]), .A3(pc[0]), .A4(n446), .Y(
        n451) );
  AND2X1_LVT U570 ( .A1(n823), .A2(inst[20]), .Y(n450) );
  AND2X1_LVT U574 ( .A1(n448), .A2(n447), .Y(br_addr[0]) );
  AO22X1_LVT U575 ( .A1(inst[3]), .A2(inst[21]), .A3(n492), .A4(inst[8]), .Y(
        n449) );
  AO21X1_LVT U576 ( .A1(n823), .A2(inst[21]), .A3(n449), .Y(n456) );
  AO22X1_LVT U578 ( .A1(n823), .A2(reg_data1[1]), .A3(pc[1]), .A4(n446), .Y(
        n455) );
  HADDX1_LVT U579 ( .A0(n451), .B0(n450), .C1(n454), .SO(n448) );
  AND2X1_LVT U580 ( .A1(n452), .A2(n447), .Y(br_addr[1]) );
  AO22X1_LVT U581 ( .A1(inst[3]), .A2(inst[22]), .A3(n492), .A4(inst[9]), .Y(
        n453) );
  AO21X1_LVT U582 ( .A1(n823), .A2(inst[22]), .A3(n453), .Y(n461) );
  AO22X1_LVT U583 ( .A1(n823), .A2(reg_data1[2]), .A3(pc[2]), .A4(n446), .Y(
        n460) );
  FADDX1_LVT U584 ( .A(n456), .B(n455), .CI(n454), .CO(n459), .S(n452) );
  AND2X1_LVT U585 ( .A1(n457), .A2(n447), .Y(br_addr[2]) );
  AO22X1_LVT U586 ( .A1(inst[3]), .A2(inst[23]), .A3(n492), .A4(inst[10]), .Y(
        n458) );
  AO21X1_LVT U587 ( .A1(n823), .A2(inst[23]), .A3(n458), .Y(n466) );
  AO22X1_LVT U589 ( .A1(n823), .A2(reg_data1[3]), .A3(n446), .A4(pc[3]), .Y(
        n465) );
  FADDX1_LVT U590 ( .A(n461), .B(n460), .CI(n459), .CO(n464), .S(n457) );
  AND2X1_LVT U591 ( .A1(n462), .A2(n447), .Y(br_addr[3]) );
  AO22X1_LVT U592 ( .A1(inst[3]), .A2(inst[24]), .A3(n492), .A4(inst[11]), .Y(
        n463) );
  AO21X1_LVT U593 ( .A1(n823), .A2(inst[24]), .A3(n463), .Y(n470) );
  AO22X1_LVT U594 ( .A1(n823), .A2(reg_data1[4]), .A3(n446), .A4(pc[4]), .Y(
        n469) );
  FADDX1_LVT U595 ( .A(n466), .B(n465), .CI(n464), .CO(n468), .S(n462) );
  AND2X1_LVT U596 ( .A1(n467), .A2(n447), .Y(br_addr[4]) );
  AO22X1_LVT U597 ( .A1(n823), .A2(reg_data1[5]), .A3(n446), .A4(pc[5]), .Y(
        n473) );
  FADDX1_LVT U598 ( .A(n470), .B(n469), .CI(n468), .CO(n472), .S(n467) );
  AND2X1_LVT U599 ( .A1(n471), .A2(n447), .Y(br_addr[5]) );
  AO22X1_LVT U600 ( .A1(n823), .A2(reg_data1[6]), .A3(n446), .A4(pc[6]), .Y(
        n476) );
  FADDX1_LVT U601 ( .A(inst[25]), .B(n473), .CI(n472), .CO(n475), .S(n471) );
  AND2X1_LVT U602 ( .A1(n474), .A2(n447), .Y(br_addr[6]) );
  AO22X1_LVT U603 ( .A1(n823), .A2(reg_data1[7]), .A3(n446), .A4(pc[7]), .Y(
        n479) );
  FADDX1_LVT U604 ( .A(inst[26]), .B(n476), .CI(n475), .CO(n478), .S(n474) );
  AND2X1_LVT U605 ( .A1(n477), .A2(n447), .Y(br_addr[7]) );
  AO22X1_LVT U606 ( .A1(n823), .A2(reg_data1[8]), .A3(n446), .A4(pc[8]), .Y(
        n482) );
  FADDX1_LVT U607 ( .A(inst[27]), .B(n479), .CI(n478), .CO(n481), .S(n477) );
  AND2X1_LVT U608 ( .A1(n480), .A2(n447), .Y(br_addr[8]) );
  AO22X1_LVT U609 ( .A1(n823), .A2(reg_data1[9]), .A3(pc[9]), .A4(n446), .Y(
        n485) );
  FADDX1_LVT U610 ( .A(inst[28]), .B(n482), .CI(n481), .CO(n484), .S(n480) );
  AND2X1_LVT U611 ( .A1(n483), .A2(n447), .Y(br_addr[9]) );
  AO22X1_LVT U612 ( .A1(n823), .A2(reg_data1[10]), .A3(pc[10]), .A4(n446), .Y(
        n490) );
  FADDX1_LVT U613 ( .A(inst[29]), .B(n485), .CI(n484), .CO(n489), .S(n483) );
  AND2X1_LVT U614 ( .A1(n486), .A2(n447), .Y(br_addr[10]) );
  NAND2X0_LVT U616 ( .A1(n822), .A2(inst[31]), .Y(n493) );
  AOI22X1_LVT U617 ( .A1(n492), .A2(inst[7]), .A3(inst[3]), .A4(inst[20]), .Y(
        n488) );
  NAND2X0_LVT U618 ( .A1(n493), .A2(n488), .Y(n497) );
  AO22X1_LVT U619 ( .A1(n823), .A2(reg_data1[11]), .A3(pc[11]), .A4(n446), .Y(
        n496) );
  FADDX1_LVT U620 ( .A(inst[30]), .B(n490), .CI(n489), .CO(n495), .S(n486) );
  AND2X1_LVT U621 ( .A1(n491), .A2(n447), .Y(br_addr[11]) );
  NAND2X0_LVT U622 ( .A1(n492), .A2(inst[31]), .Y(n494) );
  NAND2X0_LVT U623 ( .A1(n494), .A2(n493), .Y(n524) );
  AO21X1_LVT U624 ( .A1(inst[3]), .A2(inst[12]), .A3(n524), .Y(n501) );
  AO22X1_LVT U625 ( .A1(n823), .A2(reg_data1[12]), .A3(pc[12]), .A4(n446), .Y(
        n500) );
  FADDX1_LVT U626 ( .A(n497), .B(n496), .CI(n495), .CO(n499), .S(n491) );
  AND2X1_LVT U627 ( .A1(n498), .A2(n447), .Y(br_addr[12]) );
  AO21X1_LVT U628 ( .A1(inst[13]), .A2(inst[3]), .A3(n524), .Y(n505) );
  AO22X1_LVT U629 ( .A1(n823), .A2(reg_data1[13]), .A3(pc[13]), .A4(n446), .Y(
        n504) );
  FADDX1_LVT U630 ( .A(n501), .B(n500), .CI(n499), .CO(n503), .S(n498) );
  AND2X1_LVT U631 ( .A1(n502), .A2(n447), .Y(br_addr[13]) );
  AO21X1_LVT U632 ( .A1(inst[3]), .A2(N94), .A3(n524), .Y(n510) );
  AO22X1_LVT U633 ( .A1(n822), .A2(reg_data1[14]), .A3(pc[14]), .A4(n446), .Y(
        n509) );
  FADDX1_LVT U634 ( .A(n505), .B(n504), .CI(n503), .CO(n508), .S(n502) );
  AND2X1_LVT U635 ( .A1(n507), .A2(n447), .Y(br_addr[14]) );
  AO21X1_LVT U636 ( .A1(inst[3]), .A2(inst[15]), .A3(n524), .Y(n514) );
  AO22X1_LVT U637 ( .A1(n822), .A2(reg_data1[15]), .A3(pc[15]), .A4(n446), .Y(
        n513) );
  FADDX1_LVT U638 ( .A(n510), .B(n509), .CI(n508), .CO(n512), .S(n507) );
  AND2X1_LVT U640 ( .A1(n511), .A2(n447), .Y(br_addr[15]) );
  AO21X1_LVT U641 ( .A1(inst[3]), .A2(inst[16]), .A3(n524), .Y(n518) );
  AO22X1_LVT U642 ( .A1(n822), .A2(reg_data1[16]), .A3(pc[16]), .A4(n446), .Y(
        n517) );
  FADDX1_LVT U643 ( .A(n514), .B(n513), .CI(n512), .CO(n516), .S(n511) );
  AND2X1_LVT U644 ( .A1(n515), .A2(n447), .Y(br_addr[16]) );
  AO21X1_LVT U645 ( .A1(inst[3]), .A2(inst[17]), .A3(n524), .Y(n522) );
  AO22X1_LVT U646 ( .A1(n822), .A2(reg_data1[17]), .A3(pc[17]), .A4(n446), .Y(
        n521) );
  FADDX1_LVT U647 ( .A(n518), .B(n517), .CI(n516), .CO(n520), .S(n515) );
  AND2X1_LVT U648 ( .A1(n519), .A2(n447), .Y(br_addr[17]) );
  AO21X1_LVT U649 ( .A1(inst[3]), .A2(inst[18]), .A3(n524), .Y(n527) );
  AO22X1_LVT U650 ( .A1(n822), .A2(reg_data1[18]), .A3(pc[18]), .A4(n446), .Y(
        n526) );
  FADDX1_LVT U651 ( .A(n522), .B(n521), .CI(n520), .CO(n525), .S(n519) );
  AND2X1_LVT U652 ( .A1(n523), .A2(n447), .Y(br_addr[18]) );
  AO21X1_LVT U653 ( .A1(inst[3]), .A2(inst[19]), .A3(n524), .Y(n531) );
  AO22X1_LVT U654 ( .A1(n822), .A2(reg_data1[19]), .A3(pc[19]), .A4(n446), .Y(
        n530) );
  FADDX1_LVT U655 ( .A(n527), .B(n526), .CI(n525), .CO(n529), .S(n523) );
  AND2X1_LVT U656 ( .A1(n528), .A2(n447), .Y(br_addr[19]) );
  AO22X1_LVT U657 ( .A1(n822), .A2(reg_data1[20]), .A3(pc[20]), .A4(n446), .Y(
        n534) );
  FADDX1_LVT U658 ( .A(n531), .B(n530), .CI(n529), .CO(n533), .S(n528) );
  AND2X1_LVT U659 ( .A1(n532), .A2(n447), .Y(br_addr[20]) );
  AO22X1_LVT U660 ( .A1(n822), .A2(reg_data1[21]), .A3(pc[21]), .A4(n446), .Y(
        n537) );
  FADDX1_LVT U661 ( .A(n534), .B(inst[31]), .CI(n533), .CO(n536), .S(n532) );
  AND2X1_LVT U662 ( .A1(n535), .A2(n447), .Y(br_addr[21]) );
  AO22X1_LVT U663 ( .A1(n822), .A2(reg_data1[22]), .A3(pc[22]), .A4(n446), .Y(
        n540) );
  FADDX1_LVT U664 ( .A(n537), .B(inst[31]), .CI(n536), .CO(n539), .S(n535) );
  AND2X1_LVT U665 ( .A1(n538), .A2(n447), .Y(br_addr[22]) );
  AO22X1_LVT U666 ( .A1(n822), .A2(reg_data1[23]), .A3(pc[23]), .A4(n446), .Y(
        n544) );
  FADDX1_LVT U667 ( .A(n540), .B(inst[31]), .CI(n539), .CO(n543), .S(n538) );
  AND2X1_LVT U668 ( .A1(n541), .A2(n447), .Y(br_addr[23]) );
  AO22X1_LVT U669 ( .A1(n822), .A2(reg_data1[24]), .A3(pc[24]), .A4(n446), .Y(
        n547) );
  FADDX1_LVT U670 ( .A(n544), .B(inst[31]), .CI(n543), .CO(n546), .S(n541) );
  AND2X1_LVT U671 ( .A1(n545), .A2(n447), .Y(br_addr[24]) );
  AO22X1_LVT U672 ( .A1(n822), .A2(reg_data1[25]), .A3(n446), .A4(pc[25]), .Y(
        n550) );
  FADDX1_LVT U673 ( .A(n547), .B(inst[31]), .CI(n546), .CO(n549), .S(n545) );
  AND2X1_LVT U674 ( .A1(n548), .A2(n447), .Y(br_addr[25]) );
  AO22X1_LVT U675 ( .A1(n822), .A2(reg_data1[26]), .A3(n446), .A4(pc[26]), .Y(
        n553) );
  FADDX1_LVT U676 ( .A(n550), .B(inst[31]), .CI(n549), .CO(n552), .S(n548) );
  AND2X1_LVT U677 ( .A1(n551), .A2(n447), .Y(br_addr[26]) );
  AO22X1_LVT U678 ( .A1(n822), .A2(reg_data1[27]), .A3(n446), .A4(pc[27]), .Y(
        n556) );
  FADDX1_LVT U679 ( .A(n553), .B(inst[31]), .CI(n552), .CO(n555), .S(n551) );
  AND2X1_LVT U680 ( .A1(n554), .A2(n447), .Y(br_addr[27]) );
  AO22X1_LVT U681 ( .A1(n822), .A2(reg_data1[28]), .A3(n446), .A4(pc[28]), .Y(
        n561) );
  FADDX1_LVT U682 ( .A(n556), .B(inst[31]), .CI(n555), .CO(n560), .S(n554) );
  AND2X1_LVT U683 ( .A1(n557), .A2(n447), .Y(br_addr[28]) );
  AO22X1_LVT U685 ( .A1(n822), .A2(reg_data1[29]), .A3(n446), .A4(pc[29]), .Y(
        n566) );
  FADDX1_LVT U686 ( .A(n561), .B(inst[31]), .CI(n560), .CO(n565), .S(n557) );
  AND2X1_LVT U687 ( .A1(n563), .A2(n447), .Y(br_addr[29]) );
  AO22X1_LVT U688 ( .A1(n823), .A2(reg_data1[30]), .A3(n446), .A4(pc[30]), .Y(
        n570) );
  FADDX1_LVT U689 ( .A(n566), .B(inst[31]), .CI(n565), .CO(n569), .S(n563) );
  AND2X1_LVT U691 ( .A1(n568), .A2(n447), .Y(br_addr[30]) );
  FADDX1_LVT U692 ( .A(n570), .B(inst[31]), .CI(n569), .CO(n575), .S(n568) );
  AO22X1_LVT U693 ( .A1(n822), .A2(reg_data1[31]), .A3(n446), .A4(pc[31]), .Y(
        n573) );
  XOR2X1_LVT U694 ( .A1(inst[31]), .A2(n573), .Y(n574) );
  XOR2X1_LVT U695 ( .A1(n575), .A2(n574), .Y(n577) );
  AND2X1_LVT U696 ( .A1(n577), .A2(n447), .Y(br_addr[31]) );
  NAND2X0_LVT U700 ( .A1(n579), .A2(ex_we), .Y(n595) );
  AOI22X1_LVT U701 ( .A1(n582), .A2(mem_reg_waddr[2]), .A3(n581), .A4(
        mem_reg_waddr[4]), .Y(n580) );
  OA221X1_LVT U702 ( .A1(n582), .A2(mem_reg_waddr[2]), .A3(n581), .A4(
        mem_reg_waddr[4]), .A5(n580), .Y(n592) );
  OA221X1_LVT U703 ( .A1(reg_addr1[1]), .A2(n584), .A3(n583), .A4(
        mem_reg_waddr[1]), .A5(mem_we), .Y(n591) );
  OA22X1_LVT U704 ( .A1(reg_addr1[0]), .A2(n586), .A3(reg_addr1[3]), .A4(n585), 
        .Y(n587) );
  OA221X1_LVT U705 ( .A1(n589), .A2(mem_reg_waddr[0]), .A3(n588), .A4(
        mem_reg_waddr[3]), .A5(n587), .Y(n590) );
  NAND4X0_LVT U706 ( .A1(n592), .A2(n591), .A3(n590), .A4(re1), .Y(n594) );
  INVX1_LVT U710 ( .A(n594), .Y(n596) );
  AO222X1_LVT U713 ( .A1(ex_reg_wdata[0]), .A2(n578), .A3(n593), .A4(
        reg_data1[0]), .A5(mem_reg_wdata[0]), .A6(n597), .Y(N635) );
  AO222X1_LVT U716 ( .A1(n578), .A2(ex_reg_wdata[1]), .A3(n597), .A4(
        mem_reg_wdata[1]), .A5(reg_data1[1]), .A6(n593), .Y(N636) );
  AO222X1_LVT U717 ( .A1(n578), .A2(ex_reg_wdata[2]), .A3(n597), .A4(
        mem_reg_wdata[2]), .A5(reg_data1[2]), .A6(n593), .Y(N637) );
  AO222X1_LVT U718 ( .A1(n578), .A2(ex_reg_wdata[3]), .A3(n597), .A4(
        mem_reg_wdata[3]), .A5(reg_data1[3]), .A6(n593), .Y(N638) );
  AO222X1_LVT U719 ( .A1(n578), .A2(ex_reg_wdata[4]), .A3(n597), .A4(
        mem_reg_wdata[4]), .A5(reg_data1[4]), .A6(n593), .Y(N639) );
  AO222X1_LVT U720 ( .A1(n578), .A2(ex_reg_wdata[5]), .A3(n597), .A4(
        mem_reg_wdata[5]), .A5(reg_data1[5]), .A6(n593), .Y(N640) );
  AO222X1_LVT U721 ( .A1(n578), .A2(ex_reg_wdata[6]), .A3(n597), .A4(
        mem_reg_wdata[6]), .A5(reg_data1[6]), .A6(n593), .Y(N641) );
  AO222X1_LVT U722 ( .A1(n578), .A2(ex_reg_wdata[7]), .A3(n597), .A4(
        mem_reg_wdata[7]), .A5(reg_data1[7]), .A6(n593), .Y(N642) );
  AO222X1_LVT U723 ( .A1(n578), .A2(ex_reg_wdata[8]), .A3(n597), .A4(
        mem_reg_wdata[8]), .A5(reg_data1[8]), .A6(n593), .Y(N643) );
  AO222X1_LVT U724 ( .A1(n578), .A2(ex_reg_wdata[9]), .A3(n597), .A4(
        mem_reg_wdata[9]), .A5(reg_data1[9]), .A6(n593), .Y(N644) );
  AO222X1_LVT U725 ( .A1(n578), .A2(ex_reg_wdata[10]), .A3(n597), .A4(
        mem_reg_wdata[10]), .A5(reg_data1[10]), .A6(n593), .Y(N645) );
  AO222X1_LVT U726 ( .A1(n578), .A2(ex_reg_wdata[11]), .A3(n597), .A4(
        mem_reg_wdata[11]), .A5(reg_data1[11]), .A6(n593), .Y(N646) );
  AO22X1_LVT U727 ( .A1(n578), .A2(ex_reg_wdata[12]), .A3(n597), .A4(
        mem_reg_wdata[12]), .Y(n599) );
  AO22X1_LVT U728 ( .A1(inst[12]), .A2(n820), .A3(n593), .A4(reg_data1[12]), 
        .Y(n598) );
  OR2X1_LVT U729 ( .A1(n599), .A2(n598), .Y(N647) );
  AO22X1_LVT U730 ( .A1(n578), .A2(ex_reg_wdata[13]), .A3(n597), .A4(
        mem_reg_wdata[13]), .Y(n601) );
  AO22X1_LVT U731 ( .A1(inst[13]), .A2(n820), .A3(n593), .A4(reg_data1[13]), 
        .Y(n600) );
  OR2X1_LVT U732 ( .A1(n601), .A2(n600), .Y(N648) );
  AO22X1_LVT U733 ( .A1(n578), .A2(ex_reg_wdata[14]), .A3(n597), .A4(
        mem_reg_wdata[14]), .Y(n604) );
  AO22X1_LVT U734 ( .A1(N94), .A2(n820), .A3(n593), .A4(reg_data1[14]), .Y(
        n603) );
  OR2X1_LVT U735 ( .A1(n604), .A2(n603), .Y(N649) );
  AO22X1_LVT U737 ( .A1(n578), .A2(ex_reg_wdata[15]), .A3(n597), .A4(
        mem_reg_wdata[15]), .Y(n606) );
  AO22X1_LVT U738 ( .A1(inst[15]), .A2(n820), .A3(n593), .A4(reg_data1[15]), 
        .Y(n605) );
  OR2X1_LVT U739 ( .A1(n606), .A2(n605), .Y(N650) );
  AO22X1_LVT U740 ( .A1(n578), .A2(ex_reg_wdata[16]), .A3(n597), .A4(
        mem_reg_wdata[16]), .Y(n608) );
  AO22X1_LVT U741 ( .A1(inst[16]), .A2(n820), .A3(n593), .A4(reg_data1[16]), 
        .Y(n607) );
  OR2X1_LVT U742 ( .A1(n608), .A2(n607), .Y(N651) );
  AO22X1_LVT U743 ( .A1(n578), .A2(ex_reg_wdata[17]), .A3(n597), .A4(
        mem_reg_wdata[17]), .Y(n610) );
  AO22X1_LVT U744 ( .A1(inst[17]), .A2(n820), .A3(n593), .A4(reg_data1[17]), 
        .Y(n609) );
  OR2X1_LVT U745 ( .A1(n610), .A2(n609), .Y(N652) );
  AO22X1_LVT U746 ( .A1(n578), .A2(ex_reg_wdata[18]), .A3(n597), .A4(
        mem_reg_wdata[18]), .Y(n612) );
  AO22X1_LVT U747 ( .A1(inst[18]), .A2(n820), .A3(n593), .A4(reg_data1[18]), 
        .Y(n611) );
  OR2X1_LVT U748 ( .A1(n612), .A2(n611), .Y(N653) );
  AO22X1_LVT U749 ( .A1(n578), .A2(ex_reg_wdata[19]), .A3(n597), .A4(
        mem_reg_wdata[19]), .Y(n614) );
  AO22X1_LVT U750 ( .A1(inst[19]), .A2(n820), .A3(n593), .A4(reg_data1[19]), 
        .Y(n613) );
  OR2X1_LVT U751 ( .A1(n614), .A2(n613), .Y(N654) );
  AO22X1_LVT U752 ( .A1(n578), .A2(ex_reg_wdata[20]), .A3(n597), .A4(
        mem_reg_wdata[20]), .Y(n616) );
  AO22X1_LVT U753 ( .A1(n593), .A2(reg_data1[20]), .A3(n820), .A4(inst[20]), 
        .Y(n615) );
  OR2X1_LVT U754 ( .A1(n616), .A2(n615), .Y(N655) );
  AO22X1_LVT U755 ( .A1(n578), .A2(ex_reg_wdata[21]), .A3(n597), .A4(
        mem_reg_wdata[21]), .Y(n620) );
  AO22X1_LVT U757 ( .A1(n593), .A2(reg_data1[21]), .A3(n820), .A4(inst[21]), 
        .Y(n619) );
  OR2X1_LVT U758 ( .A1(n620), .A2(n619), .Y(N656) );
  AO22X1_LVT U759 ( .A1(n578), .A2(ex_reg_wdata[22]), .A3(n597), .A4(
        mem_reg_wdata[22]), .Y(n622) );
  AO22X1_LVT U760 ( .A1(n593), .A2(reg_data1[22]), .A3(n820), .A4(inst[22]), 
        .Y(n621) );
  OR2X1_LVT U761 ( .A1(n622), .A2(n621), .Y(N657) );
  AO22X1_LVT U762 ( .A1(n578), .A2(ex_reg_wdata[23]), .A3(n597), .A4(
        mem_reg_wdata[23]), .Y(n624) );
  AO22X1_LVT U763 ( .A1(n593), .A2(reg_data1[23]), .A3(n820), .A4(inst[23]), 
        .Y(n623) );
  OR2X1_LVT U764 ( .A1(n624), .A2(n623), .Y(N658) );
  AO22X1_LVT U765 ( .A1(n578), .A2(ex_reg_wdata[24]), .A3(n597), .A4(
        mem_reg_wdata[24]), .Y(n626) );
  AO22X1_LVT U766 ( .A1(n593), .A2(reg_data1[24]), .A3(n820), .A4(inst[24]), 
        .Y(n625) );
  OR2X1_LVT U767 ( .A1(n626), .A2(n625), .Y(N659) );
  AO22X1_LVT U768 ( .A1(n578), .A2(ex_reg_wdata[25]), .A3(n597), .A4(
        mem_reg_wdata[25]), .Y(n628) );
  AO22X1_LVT U769 ( .A1(inst[25]), .A2(n820), .A3(n593), .A4(reg_data1[25]), 
        .Y(n627) );
  OR2X1_LVT U770 ( .A1(n628), .A2(n627), .Y(N660) );
  AO22X1_LVT U771 ( .A1(n578), .A2(ex_reg_wdata[26]), .A3(n597), .A4(
        mem_reg_wdata[26]), .Y(n630) );
  AO22X1_LVT U772 ( .A1(inst[26]), .A2(n820), .A3(n593), .A4(reg_data1[26]), 
        .Y(n629) );
  OR2X1_LVT U773 ( .A1(n630), .A2(n629), .Y(N661) );
  AO22X1_LVT U774 ( .A1(n578), .A2(ex_reg_wdata[27]), .A3(n597), .A4(
        mem_reg_wdata[27]), .Y(n632) );
  AO22X1_LVT U775 ( .A1(inst[27]), .A2(n820), .A3(n593), .A4(reg_data1[27]), 
        .Y(n631) );
  OR2X1_LVT U776 ( .A1(n632), .A2(n631), .Y(N662) );
  AO22X1_LVT U777 ( .A1(n578), .A2(ex_reg_wdata[28]), .A3(n597), .A4(
        mem_reg_wdata[28]), .Y(n634) );
  AO22X1_LVT U778 ( .A1(inst[28]), .A2(n820), .A3(n593), .A4(reg_data1[28]), 
        .Y(n633) );
  OR2X1_LVT U779 ( .A1(n634), .A2(n633), .Y(N663) );
  AO22X1_LVT U780 ( .A1(n578), .A2(ex_reg_wdata[29]), .A3(n597), .A4(
        mem_reg_wdata[29]), .Y(n636) );
  AO22X1_LVT U781 ( .A1(inst[29]), .A2(n820), .A3(n593), .A4(reg_data1[29]), 
        .Y(n635) );
  OR2X1_LVT U782 ( .A1(n636), .A2(n635), .Y(N664) );
  AO22X1_LVT U783 ( .A1(n578), .A2(ex_reg_wdata[30]), .A3(n597), .A4(
        mem_reg_wdata[30]), .Y(n641) );
  AO22X1_LVT U784 ( .A1(n593), .A2(reg_data1[30]), .A3(n820), .A4(inst[30]), 
        .Y(n640) );
  OR2X1_LVT U785 ( .A1(n641), .A2(n640), .Y(N665) );
  AO22X1_LVT U787 ( .A1(n578), .A2(ex_reg_wdata[31]), .A3(n597), .A4(
        mem_reg_wdata[31]), .Y(n648) );
  AO22X1_LVT U788 ( .A1(inst[31]), .A2(n820), .A3(n593), .A4(reg_data1[31]), 
        .Y(n647) );
  OR2X1_LVT U789 ( .A1(n648), .A2(n647), .Y(N666) );
  AOI22X1_LVT U790 ( .A1(mem_reg_wdata[12]), .A2(n274), .A3(ex_reg_wdata[12]), 
        .A4(n257), .Y(n651) );
  NAND2X0_LVT U791 ( .A1(n267), .A2(reg_data2[12]), .Y(n650) );
  NAND2X0_LVT U793 ( .A1(pc[12]), .A2(n665), .Y(n649) );
  NAND4X0_LVT U794 ( .A1(n651), .A2(n650), .A3(n839), .A4(n649), .Y(N708) );
  AOI22X1_LVT U796 ( .A1(mem_reg_wdata[13]), .A2(n274), .A3(ex_reg_wdata[13]), 
        .A4(n257), .Y(n655) );
  NAND2X0_LVT U798 ( .A1(n267), .A2(reg_data2[13]), .Y(n654) );
  NAND2X0_LVT U799 ( .A1(pc[13]), .A2(n665), .Y(n653) );
  NAND4X0_LVT U800 ( .A1(n655), .A2(n839), .A3(n654), .A4(n653), .Y(N709) );
  AOI22X1_LVT U801 ( .A1(mem_reg_wdata[14]), .A2(n274), .A3(ex_reg_wdata[14]), 
        .A4(n257), .Y(n659) );
  NAND2X0_LVT U803 ( .A1(n267), .A2(reg_data2[14]), .Y(n658) );
  NAND2X0_LVT U804 ( .A1(pc[14]), .A2(n665), .Y(n657) );
  NAND4X0_LVT U805 ( .A1(n659), .A2(n839), .A3(n658), .A4(n657), .Y(N710) );
  AOI22X1_LVT U806 ( .A1(mem_reg_wdata[15]), .A2(n274), .A3(ex_reg_wdata[15]), 
        .A4(n257), .Y(n663) );
  NAND2X0_LVT U807 ( .A1(n267), .A2(reg_data2[15]), .Y(n662) );
  NAND2X0_LVT U808 ( .A1(pc[15]), .A2(n665), .Y(n661) );
  NAND4X0_LVT U809 ( .A1(n663), .A2(n839), .A3(n662), .A4(n661), .Y(N711) );
  AOI22X1_LVT U811 ( .A1(mem_reg_wdata[16]), .A2(n274), .A3(ex_reg_wdata[16]), 
        .A4(n257), .Y(n668) );
  NAND2X0_LVT U812 ( .A1(n267), .A2(reg_data2[16]), .Y(n667) );
  NAND2X0_LVT U814 ( .A1(pc[16]), .A2(n665), .Y(n666) );
  NAND4X0_LVT U815 ( .A1(n668), .A2(n839), .A3(n667), .A4(n666), .Y(N712) );
  AOI22X1_LVT U816 ( .A1(mem_reg_wdata[17]), .A2(n274), .A3(ex_reg_wdata[17]), 
        .A4(n257), .Y(n671) );
  NAND2X0_LVT U817 ( .A1(n267), .A2(reg_data2[17]), .Y(n670) );
  NAND2X0_LVT U818 ( .A1(pc[17]), .A2(n665), .Y(n669) );
  NAND4X0_LVT U819 ( .A1(n671), .A2(n839), .A3(n670), .A4(n669), .Y(N713) );
  AOI22X1_LVT U820 ( .A1(mem_reg_wdata[18]), .A2(n274), .A3(ex_reg_wdata[18]), 
        .A4(n257), .Y(n674) );
  NAND2X0_LVT U821 ( .A1(n267), .A2(reg_data2[18]), .Y(n673) );
  NAND2X0_LVT U822 ( .A1(pc[18]), .A2(n665), .Y(n672) );
  NAND4X0_LVT U823 ( .A1(n674), .A2(n839), .A3(n673), .A4(n672), .Y(N714) );
  AOI22X1_LVT U824 ( .A1(mem_reg_wdata[19]), .A2(n274), .A3(ex_reg_wdata[19]), 
        .A4(n257), .Y(n677) );
  NAND2X0_LVT U825 ( .A1(n267), .A2(reg_data2[19]), .Y(n676) );
  NAND2X0_LVT U826 ( .A1(pc[19]), .A2(n665), .Y(n675) );
  NAND4X0_LVT U827 ( .A1(n677), .A2(n839), .A3(n676), .A4(n675), .Y(N715) );
  AOI22X1_LVT U828 ( .A1(mem_reg_wdata[20]), .A2(n274), .A3(ex_reg_wdata[20]), 
        .A4(n257), .Y(n680) );
  NAND2X0_LVT U829 ( .A1(n267), .A2(reg_data2[20]), .Y(n679) );
  NAND2X0_LVT U830 ( .A1(pc[20]), .A2(n665), .Y(n678) );
  NAND4X0_LVT U831 ( .A1(n680), .A2(n839), .A3(n679), .A4(n678), .Y(N716) );
  AOI22X1_LVT U832 ( .A1(mem_reg_wdata[21]), .A2(n274), .A3(ex_reg_wdata[21]), 
        .A4(n257), .Y(n683) );
  NAND2X0_LVT U833 ( .A1(n267), .A2(reg_data2[21]), .Y(n682) );
  NAND2X0_LVT U834 ( .A1(pc[21]), .A2(n665), .Y(n681) );
  NAND4X0_LVT U835 ( .A1(n683), .A2(n839), .A3(n682), .A4(n681), .Y(N717) );
  AOI22X1_LVT U836 ( .A1(mem_reg_wdata[22]), .A2(n274), .A3(ex_reg_wdata[22]), 
        .A4(n257), .Y(n686) );
  NAND2X0_LVT U837 ( .A1(n267), .A2(reg_data2[22]), .Y(n685) );
  NAND2X0_LVT U838 ( .A1(pc[22]), .A2(n665), .Y(n684) );
  NAND4X0_LVT U839 ( .A1(n686), .A2(n839), .A3(n685), .A4(n684), .Y(N718) );
  AOI22X1_LVT U840 ( .A1(mem_reg_wdata[23]), .A2(n274), .A3(ex_reg_wdata[23]), 
        .A4(n257), .Y(n689) );
  NAND2X0_LVT U841 ( .A1(n267), .A2(reg_data2[23]), .Y(n688) );
  NAND2X0_LVT U842 ( .A1(pc[23]), .A2(n665), .Y(n687) );
  NAND4X0_LVT U843 ( .A1(n689), .A2(n839), .A3(n688), .A4(n687), .Y(N719) );
  AOI22X1_LVT U844 ( .A1(mem_reg_wdata[24]), .A2(n274), .A3(ex_reg_wdata[24]), 
        .A4(n257), .Y(n692) );
  NAND2X0_LVT U845 ( .A1(n267), .A2(reg_data2[24]), .Y(n691) );
  NAND2X0_LVT U846 ( .A1(pc[24]), .A2(n665), .Y(n690) );
  NAND4X0_LVT U847 ( .A1(n692), .A2(n839), .A3(n691), .A4(n690), .Y(N720) );
  AOI22X1_LVT U848 ( .A1(mem_reg_wdata[25]), .A2(n274), .A3(ex_reg_wdata[25]), 
        .A4(n257), .Y(n695) );
  NAND2X0_LVT U849 ( .A1(n267), .A2(reg_data2[25]), .Y(n694) );
  NAND2X0_LVT U850 ( .A1(pc[25]), .A2(n665), .Y(n693) );
  NAND4X0_LVT U851 ( .A1(n695), .A2(n839), .A3(n694), .A4(n693), .Y(N721) );
  AOI22X1_LVT U852 ( .A1(mem_reg_wdata[26]), .A2(n274), .A3(ex_reg_wdata[26]), 
        .A4(n257), .Y(n698) );
  NAND2X0_LVT U853 ( .A1(n267), .A2(reg_data2[26]), .Y(n697) );
  NAND2X0_LVT U854 ( .A1(pc[26]), .A2(n665), .Y(n696) );
  NAND4X0_LVT U855 ( .A1(n698), .A2(n722), .A3(n697), .A4(n696), .Y(N722) );
  AOI22X1_LVT U856 ( .A1(mem_reg_wdata[27]), .A2(n274), .A3(ex_reg_wdata[27]), 
        .A4(n257), .Y(n701) );
  NAND2X0_LVT U857 ( .A1(n267), .A2(reg_data2[27]), .Y(n700) );
  NAND2X0_LVT U858 ( .A1(pc[27]), .A2(n665), .Y(n699) );
  NAND4X0_LVT U859 ( .A1(n701), .A2(n722), .A3(n700), .A4(n699), .Y(N723) );
  AOI22X1_LVT U860 ( .A1(mem_reg_wdata[28]), .A2(n274), .A3(ex_reg_wdata[28]), 
        .A4(n257), .Y(n705) );
  NAND2X0_LVT U861 ( .A1(n267), .A2(reg_data2[28]), .Y(n704) );
  NAND2X0_LVT U862 ( .A1(pc[28]), .A2(n665), .Y(n703) );
  NAND4X0_LVT U863 ( .A1(n705), .A2(n722), .A3(n704), .A4(n703), .Y(N724) );
  AOI22X1_LVT U864 ( .A1(mem_reg_wdata[29]), .A2(n274), .A3(ex_reg_wdata[29]), 
        .A4(n257), .Y(n709) );
  NAND2X0_LVT U865 ( .A1(n267), .A2(reg_data2[29]), .Y(n708) );
  NAND2X0_LVT U866 ( .A1(pc[29]), .A2(n665), .Y(n707) );
  NAND4X0_LVT U867 ( .A1(n709), .A2(n722), .A3(n708), .A4(n707), .Y(N725) );
  AOI22X1_LVT U868 ( .A1(mem_reg_wdata[30]), .A2(n274), .A3(ex_reg_wdata[30]), 
        .A4(n257), .Y(n714) );
  NAND2X0_LVT U869 ( .A1(n267), .A2(reg_data2[30]), .Y(n713) );
  NAND2X0_LVT U870 ( .A1(pc[30]), .A2(n665), .Y(n712) );
  NAND4X0_LVT U871 ( .A1(n714), .A2(n722), .A3(n713), .A4(n712), .Y(N726) );
  AOI22X1_LVT U872 ( .A1(ex_reg_wdata[31]), .A2(n257), .A3(n267), .A4(
        reg_data2[31]), .Y(n723) );
  NAND2X0_LVT U874 ( .A1(mem_reg_wdata[31]), .A2(n274), .Y(n721) );
  NAND2X0_LVT U875 ( .A1(pc[31]), .A2(n665), .Y(n720) );
  NAND4X0_LVT U876 ( .A1(n723), .A2(n722), .A3(n721), .A4(n720), .Y(N727) );
  AND2X1_LVT U877 ( .A1(n821), .A2(pc[0]), .Y(link_addr[0]) );
  AND2X1_LVT U878 ( .A1(n821), .A2(pc[1]), .Y(link_addr[1]) );
  AND2X1_LVT U880 ( .A1(n821), .A2(n816), .Y(link_addr[2]) );
  OA221X1_LVT U882 ( .A1(pc[2]), .A2(pc[3]), .A3(n816), .A4(n817), .A5(n821), 
        .Y(link_addr[3]) );
  INVX1_LVT U883 ( .A(n728), .Y(n730) );
  OA221X1_LVT U885 ( .A1(pc[31]), .A2(n730), .A3(n819), .A4(n728), .A5(n821), 
        .Y(link_addr[31]) );
  INVX1_LVT U886 ( .A(n799), .Y(n732) );
  INVX1_LVT U887 ( .A(n731), .Y(n792) );
  AO22X1_LVT U888 ( .A1(n732), .A2(inst[7]), .A3(n792), .A4(inst[20]), .Y(
        mem_offset[0]) );
  AO22X1_LVT U889 ( .A1(n732), .A2(inst[8]), .A3(n792), .A4(inst[21]), .Y(
        mem_offset[1]) );
  AO22X1_LVT U890 ( .A1(n732), .A2(inst[9]), .A3(n792), .A4(inst[22]), .Y(
        mem_offset[2]) );
  AO22X1_LVT U891 ( .A1(n732), .A2(inst[10]), .A3(n792), .A4(inst[23]), .Y(
        mem_offset[3]) );
  AO22X1_LVT U892 ( .A1(n732), .A2(inst[11]), .A3(n792), .A4(inst[24]), .Y(
        mem_offset[4]) );
  AND2X1_LVT U893 ( .A1(inst[25]), .A2(n801), .Y(mem_offset[5]) );
  AND2X1_LVT U894 ( .A1(inst[26]), .A2(n801), .Y(mem_offset[6]) );
  AND2X1_LVT U895 ( .A1(inst[27]), .A2(n801), .Y(mem_offset[7]) );
  AND2X1_LVT U896 ( .A1(inst[28]), .A2(n801), .Y(mem_offset[8]) );
  AND2X1_LVT U897 ( .A1(inst[29]), .A2(n801), .Y(mem_offset[9]) );
  AND2X1_LVT U898 ( .A1(inst[30]), .A2(n801), .Y(mem_offset[10]) );
  INVX1_LVT U899 ( .A(n733), .Y(n741) );
  AO21X1_LVT U900 ( .A1(inst[2]), .A2(n748), .A3(n746), .Y(n734) );
  NAND2X0_LVT U901 ( .A1(n735), .A2(n734), .Y(n736) );
  NAND4X0_LVT U902 ( .A1(n741), .A2(n809), .A3(n740), .A4(n736), .Y(n738) );
  AND2X1_LVT U903 ( .A1(inst[7]), .A2(n738), .Y(reg_waddr[0]) );
  AND2X1_LVT U904 ( .A1(inst[8]), .A2(n738), .Y(reg_waddr[1]) );
  AND2X1_LVT U905 ( .A1(inst[9]), .A2(n738), .Y(reg_waddr[2]) );
  AND2X1_LVT U906 ( .A1(inst[10]), .A2(n738), .Y(reg_waddr[3]) );
  AND2X1_LVT U907 ( .A1(inst[11]), .A2(n738), .Y(reg_waddr[4]) );
  NAND4X0_LVT U908 ( .A1(n741), .A2(n743), .A3(n740), .A4(n739), .Y(we) );
  NAND3X0_LVT U909 ( .A1(n765), .A2(N94), .A3(n759), .Y(n742) );
  NAND2X0_LVT U910 ( .A1(n752), .A2(n742), .Y(alusel[0]) );
  AND2X1_LVT U911 ( .A1(N94), .A2(n758), .Y(n775) );
  AO222X1_LVT U912 ( .A1(n743), .A2(n775), .A3(n743), .A4(n779), .A5(n743), 
        .A6(n759), .Y(n794) );
  NAND3X0_LVT U913 ( .A1(n794), .A2(n755), .A3(n752), .Y(alusel[1]) );
  OAI21X1_LVT U914 ( .A1(n745), .A2(n758), .A3(n744), .Y(n747) );
  AO221X1_LVT U915 ( .A1(n748), .A2(inst[2]), .A3(n748), .A4(n747), .A5(n746), 
        .Y(n750) );
  AOI22X1_LVT U916 ( .A1(n751), .A2(n750), .A3(n749), .A4(n812), .Y(n800) );
  NAND3X0_LVT U917 ( .A1(n800), .A2(n755), .A3(n752), .Y(alusel[2]) );
  AOI21X1_LVT U918 ( .A1(n754), .A2(n813), .A3(n823), .Y(n757) );
  OA22X1_LVT U919 ( .A1(n757), .A2(n756), .A3(n813), .A4(n755), .Y(n773) );
  INVX1_LVT U920 ( .A(n758), .Y(n766) );
  INVX1_LVT U921 ( .A(n759), .Y(n795) );
  NAND4X0_LVT U922 ( .A1(n766), .A2(n795), .A3(n765), .A4(inst[30]), .Y(n772)
         );
  INVX1_LVT U923 ( .A(n760), .Y(n763) );
  NAND2X0_LVT U925 ( .A1(n779), .A2(n782), .Y(n761) );
  NAND3X0_LVT U926 ( .A1(n763), .A2(n836), .A3(n761), .Y(n771) );
  INVX1_LVT U927 ( .A(n764), .Y(n769) );
  INVX1_LVT U928 ( .A(n779), .Y(n768) );
  NAND4X0_LVT U929 ( .A1(inst[5]), .A2(n766), .A3(n765), .A4(inst[30]), .Y(
        n784) );
  NAND2X0_LVT U930 ( .A1(n784), .A2(n836), .Y(n767) );
  NAND3X0_LVT U931 ( .A1(n769), .A2(n768), .A3(n767), .Y(n770) );
  NAND4X0_LVT U932 ( .A1(n773), .A2(n772), .A3(n771), .A4(n770), .Y(aluop[0])
         );
  OA21X1_LVT U933 ( .A1(n836), .A2(n812), .A3(n774), .Y(n781) );
  INVX1_LVT U934 ( .A(n776), .Y(n777) );
  AO222X1_LVT U935 ( .A1(N94), .A2(n777), .A3(n812), .A4(n776), .A5(inst[12]), 
        .A6(n775), .Y(n778) );
  OA22X1_LVT U936 ( .A1(n781), .A2(n780), .A3(n779), .A4(n778), .Y(n788) );
  INVX1_LVT U937 ( .A(n781), .Y(n783) );
  OA22X1_LVT U938 ( .A1(inst[13]), .A2(n784), .A3(n783), .A4(n782), .Y(n785)
         );
  OA222X1_LVT U939 ( .A1(n799), .A2(n836), .A3(n799), .A4(n813), .A5(inst[12]), 
        .A6(n785), .Y(n787) );
  NAND2X0_LVT U940 ( .A1(n788), .A2(n787), .Y(aluop[1]) );
  NAND3X0_LVT U941 ( .A1(n802), .A2(n812), .A3(n836), .Y(n798) );
  NAND2X0_LVT U942 ( .A1(N94), .A2(inst[12]), .Y(n791) );
  NAND2X0_LVT U943 ( .A1(n792), .A2(n791), .Y(n793) );
  NAND3X0_LVT U944 ( .A1(n794), .A2(n798), .A3(n793), .Y(aluop[2]) );
  NAND3X0_LVT U945 ( .A1(N94), .A2(n796), .A3(n795), .Y(n797) );
  NAND4X0_LVT U946 ( .A1(n800), .A2(n799), .A3(n798), .A4(n797), .Y(aluop[3])
         );
  AO21X1_LVT U947 ( .A1(N94), .A2(n802), .A3(n801), .Y(aluop[4]) );
  NAND2X2_LVT U285 ( .A1(n743), .A2(n226), .Y(br) );
  AND3X4_LVT U697 ( .A1(n579), .A2(ex_we), .A3(n237), .Y(n578) );
  AND3X4_LVT U711 ( .A1(n596), .A2(n237), .A3(n595), .Y(n597) );
  AND4X4_LVT U707 ( .A1(re1), .A2(n237), .A3(n595), .A4(n594), .Y(n593) );
  AND4X4_LVT U339 ( .A1(re2), .A2(n254), .A3(n272), .A4(n271), .Y(n267) );
  AND2X4_LVT U307 ( .A1(inst[31]), .A2(n801), .Y(mem_offset[31]) );
  NAND2X4_LVT U571 ( .A1(n743), .A2(n755), .Y(n447) );
  AND2X4_LVT U346 ( .A1(n820), .A2(n269), .Y(n665) );
  NAND2X4_LVT U566 ( .A1(n445), .A2(n811), .Y(n446) );
  INVX1_LVT U3 ( .A(rst), .Y(n809) );
  INVX1_LVT U7 ( .A(ex_aluop[2]), .Y(n810) );
  INVX1_LVT U12 ( .A(inst[3]), .Y(n811) );
  INVX1_LVT U15 ( .A(N94), .Y(n812) );
  INVX1_LVT U16 ( .A(inst[12]), .Y(n813) );
  INVX1_LVT U24 ( .A(inst[13]), .Y(n814) );
  INVX1_LVT U35 ( .A(inst[21]), .Y(n815) );
  INVX1_LVT U37 ( .A(pc[2]), .Y(n816) );
  INVX1_LVT U57 ( .A(pc[3]), .Y(n817) );
  INVX1_LVT U58 ( .A(inst[24]), .Y(n818) );
  INVX1_LVT U64 ( .A(pc[31]), .Y(n819) );
  INVX2_LVT U66 ( .A(n739), .Y(n820) );
  INVX4_LVT U72 ( .A(n743), .Y(n821) );
  NBUFFX4_LVT U81 ( .A(n10), .Y(n822) );
  NBUFFX4_LVT U84 ( .A(n10), .Y(n823) );
  INVX2_LVT U142 ( .A(n246), .Y(reg_addr2[3]) );
  INVX1_LVT U161 ( .A(n582), .Y(reg_addr1[2]) );
  INVX1_LVT U290 ( .A(n588), .Y(reg_addr1[3]) );
  INVX1_LVT U300 ( .A(n581), .Y(reg_addr1[4]) );
  INVX1_LVT U301 ( .A(opv1[16]), .Y(n829) );
  INVX1_LVT U310 ( .A(opv1[17]), .Y(n830) );
  INVX1_LVT U317 ( .A(opv1[22]), .Y(n831) );
  INVX1_LVT U318 ( .A(opv1[24]), .Y(n832) );
  INVX1_LVT U320 ( .A(opv1[25]), .Y(n833) );
  AND3X4_LVT U324 ( .A1(n258), .A2(ex_we), .A3(n838), .Y(n257) );
  AND3X4_LVT U353 ( .A1(n273), .A2(n838), .A3(n272), .Y(n274) );
  NAND2X4_LVT U73 ( .A1(n751), .A2(n746), .Y(n743) );
  LATCHX2_LVT \opv1_reg[17]  ( .CLK(n835), .D(N652), .Q(opv1[17]) );
  NAND2X4_LVT U316 ( .A1(n253), .A2(n258), .Y(n254) );
  INVX2_LVT U306 ( .A(n752), .Y(n801) );
  LATCHX2_LVT \opv1_reg[16]  ( .CLK(n835), .D(N651), .Q(opv1[16]) );
  INVX2_LVT U156 ( .A(n260), .Y(reg_addr2[2]) );
  LATCHX2_LVT \opv1_reg[25]  ( .CLK(n835), .D(N660), .Q(opv1[25]) );
  NAND3X0_LVT U792 ( .A1(inst[31]), .A2(n749), .A3(n812), .Y(n722) );
  NAND2X2_LVT U299 ( .A1(n253), .A2(n579), .Y(n237) );
  NBUFFX4_LVT U321 ( .A(n814), .Y(n836) );
  NBUFFX4_LVT U322 ( .A(pc[10]), .Y(n834) );
  NBUFFX4_LVT U323 ( .A(mem_offset[31]), .Y(\mem_offset[11] ) );
  NBUFFX4_LVT U325 ( .A(n722), .Y(n839) );
  NBUFFX4_LVT U326 ( .A(n237), .Y(n835) );
  NBUFFX4_LVT U331 ( .A(n254), .Y(n838) );
endmodule


module regfile ( clk, rst, we, waddr, wdata, re1, raddr1, rdata1, re2, raddr2, 
        rdata2 );
  input [4:0] waddr;
  input [31:0] wdata;
  input [4:0] raddr1;
  output [31:0] rdata1;
  input [4:0] raddr2;
  output [31:0] rdata2;
  input clk, rst, we, re1, re2;
  wire   \regs[1][31] , \regs[1][30] , \regs[1][29] , \regs[1][28] ,
         \regs[1][27] , \regs[1][26] , \regs[1][25] , \regs[1][24] ,
         \regs[1][23] , \regs[1][22] , \regs[1][21] , \regs[1][20] ,
         \regs[1][19] , \regs[1][18] , \regs[1][17] , \regs[1][16] ,
         \regs[1][15] , \regs[1][14] , \regs[1][13] , \regs[1][12] ,
         \regs[1][11] , \regs[1][10] , \regs[1][9] , \regs[1][8] ,
         \regs[1][7] , \regs[1][6] , \regs[1][5] , \regs[1][4] , \regs[1][3] ,
         \regs[1][2] , \regs[1][1] , \regs[1][0] , \regs[2][31] ,
         \regs[2][30] , \regs[2][29] , \regs[2][28] , \regs[2][27] ,
         \regs[2][26] , \regs[2][25] , \regs[2][24] , \regs[2][23] ,
         \regs[2][22] , \regs[2][21] , \regs[2][20] , \regs[2][19] ,
         \regs[2][18] , \regs[2][17] , \regs[2][16] , \regs[2][15] ,
         \regs[2][14] , \regs[2][13] , \regs[2][12] , \regs[2][11] ,
         \regs[2][10] , \regs[2][9] , \regs[2][8] , \regs[2][7] , \regs[2][6] ,
         \regs[2][5] , \regs[2][4] , \regs[2][3] , \regs[2][2] , \regs[2][1] ,
         \regs[2][0] , \regs[3][31] , \regs[3][30] , \regs[3][29] ,
         \regs[3][28] , \regs[3][27] , \regs[3][26] , \regs[3][25] ,
         \regs[3][24] , \regs[3][23] , \regs[3][22] , \regs[3][21] ,
         \regs[3][20] , \regs[3][19] , \regs[3][18] , \regs[3][17] ,
         \regs[3][16] , \regs[3][15] , \regs[3][14] , \regs[3][13] ,
         \regs[3][12] , \regs[3][11] , \regs[3][10] , \regs[3][9] ,
         \regs[3][8] , \regs[3][7] , \regs[3][6] , \regs[3][5] , \regs[3][4] ,
         \regs[3][3] , \regs[3][2] , \regs[3][1] , \regs[3][0] , \regs[4][31] ,
         \regs[4][30] , \regs[4][29] , \regs[4][28] , \regs[4][27] ,
         \regs[4][26] , \regs[4][25] , \regs[4][24] , \regs[4][23] ,
         \regs[4][22] , \regs[4][21] , \regs[4][20] , \regs[4][19] ,
         \regs[4][18] , \regs[4][17] , \regs[4][16] , \regs[4][15] ,
         \regs[4][14] , \regs[4][13] , \regs[4][12] , \regs[4][11] ,
         \regs[4][10] , \regs[4][9] , \regs[4][8] , \regs[4][7] , \regs[4][6] ,
         \regs[4][5] , \regs[4][4] , \regs[4][3] , \regs[4][2] , \regs[4][1] ,
         \regs[4][0] , \regs[5][31] , \regs[5][30] , \regs[5][29] ,
         \regs[5][28] , \regs[5][27] , \regs[5][26] , \regs[5][25] ,
         \regs[5][24] , \regs[5][23] , \regs[5][22] , \regs[5][21] ,
         \regs[5][20] , \regs[5][19] , \regs[5][18] , \regs[5][17] ,
         \regs[5][16] , \regs[5][15] , \regs[5][14] , \regs[5][13] ,
         \regs[5][12] , \regs[5][11] , \regs[5][10] , \regs[5][9] ,
         \regs[5][8] , \regs[5][7] , \regs[5][6] , \regs[5][5] , \regs[5][4] ,
         \regs[5][3] , \regs[5][2] , \regs[5][1] , \regs[5][0] , \regs[6][31] ,
         \regs[6][30] , \regs[6][29] , \regs[6][28] , \regs[6][27] ,
         \regs[6][26] , \regs[6][25] , \regs[6][24] , \regs[6][23] ,
         \regs[6][22] , \regs[6][21] , \regs[6][20] , \regs[6][19] ,
         \regs[6][18] , \regs[6][17] , \regs[6][16] , \regs[6][15] ,
         \regs[6][14] , \regs[6][13] , \regs[6][12] , \regs[6][11] ,
         \regs[6][10] , \regs[6][9] , \regs[6][8] , \regs[6][7] , \regs[6][6] ,
         \regs[6][5] , \regs[6][4] , \regs[6][3] , \regs[6][2] , \regs[6][1] ,
         \regs[6][0] , \regs[7][31] , \regs[7][30] , \regs[7][29] ,
         \regs[7][28] , \regs[7][27] , \regs[7][26] , \regs[7][25] ,
         \regs[7][24] , \regs[7][23] , \regs[7][22] , \regs[7][21] ,
         \regs[7][20] , \regs[7][19] , \regs[7][18] , \regs[7][17] ,
         \regs[7][16] , \regs[7][15] , \regs[7][14] , \regs[7][13] ,
         \regs[7][12] , \regs[7][11] , \regs[7][10] , \regs[7][9] ,
         \regs[7][8] , \regs[7][7] , \regs[7][6] , \regs[7][5] , \regs[7][4] ,
         \regs[7][3] , \regs[7][2] , \regs[7][1] , \regs[7][0] , \regs[8][31] ,
         \regs[8][30] , \regs[8][29] , \regs[8][28] , \regs[8][27] ,
         \regs[8][26] , \regs[8][25] , \regs[8][24] , \regs[8][23] ,
         \regs[8][22] , \regs[8][21] , \regs[8][20] , \regs[8][19] ,
         \regs[8][18] , \regs[8][17] , \regs[8][16] , \regs[8][15] ,
         \regs[8][14] , \regs[8][13] , \regs[8][12] , \regs[8][11] ,
         \regs[8][10] , \regs[8][9] , \regs[8][8] , \regs[8][7] , \regs[8][6] ,
         \regs[8][5] , \regs[8][4] , \regs[8][3] , \regs[8][2] , \regs[8][1] ,
         \regs[8][0] , \regs[9][31] , \regs[9][30] , \regs[9][29] ,
         \regs[9][28] , \regs[9][27] , \regs[9][26] , \regs[9][25] ,
         \regs[9][24] , \regs[9][23] , \regs[9][22] , \regs[9][21] ,
         \regs[9][20] , \regs[9][19] , \regs[9][18] , \regs[9][17] ,
         \regs[9][16] , \regs[9][15] , \regs[9][14] , \regs[9][13] ,
         \regs[9][12] , \regs[9][11] , \regs[9][10] , \regs[9][9] ,
         \regs[9][8] , \regs[9][7] , \regs[9][6] , \regs[9][5] , \regs[9][4] ,
         \regs[9][3] , \regs[9][2] , \regs[9][1] , \regs[9][0] ,
         \regs[10][31] , \regs[10][30] , \regs[10][29] , \regs[10][28] ,
         \regs[10][27] , \regs[10][26] , \regs[10][25] , \regs[10][24] ,
         \regs[10][23] , \regs[10][22] , \regs[10][21] , \regs[10][20] ,
         \regs[10][19] , \regs[10][18] , \regs[10][17] , \regs[10][16] ,
         \regs[10][15] , \regs[10][14] , \regs[10][13] , \regs[10][12] ,
         \regs[10][11] , \regs[10][10] , \regs[10][9] , \regs[10][8] ,
         \regs[10][7] , \regs[10][6] , \regs[10][5] , \regs[10][4] ,
         \regs[10][3] , \regs[10][2] , \regs[10][1] , \regs[10][0] ,
         \regs[11][31] , \regs[11][30] , \regs[11][29] , \regs[11][28] ,
         \regs[11][27] , \regs[11][26] , \regs[11][25] , \regs[11][24] ,
         \regs[11][23] , \regs[11][22] , \regs[11][21] , \regs[11][20] ,
         \regs[11][19] , \regs[11][18] , \regs[11][17] , \regs[11][16] ,
         \regs[11][15] , \regs[11][14] , \regs[11][13] , \regs[11][12] ,
         \regs[11][11] , \regs[11][10] , \regs[11][9] , \regs[11][8] ,
         \regs[11][7] , \regs[11][6] , \regs[11][5] , \regs[11][4] ,
         \regs[11][3] , \regs[11][2] , \regs[11][1] , \regs[11][0] ,
         \regs[12][31] , \regs[12][30] , \regs[12][29] , \regs[12][28] ,
         \regs[12][27] , \regs[12][26] , \regs[12][25] , \regs[12][24] ,
         \regs[12][23] , \regs[12][22] , \regs[12][21] , \regs[12][20] ,
         \regs[12][19] , \regs[12][18] , \regs[12][17] , \regs[12][16] ,
         \regs[12][15] , \regs[12][14] , \regs[12][13] , \regs[12][12] ,
         \regs[12][11] , \regs[12][10] , \regs[12][9] , \regs[12][8] ,
         \regs[12][7] , \regs[12][6] , \regs[12][5] , \regs[12][4] ,
         \regs[12][3] , \regs[12][2] , \regs[12][1] , \regs[12][0] ,
         \regs[13][31] , \regs[13][30] , \regs[13][29] , \regs[13][28] ,
         \regs[13][27] , \regs[13][26] , \regs[13][25] , \regs[13][24] ,
         \regs[13][23] , \regs[13][22] , \regs[13][21] , \regs[13][20] ,
         \regs[13][19] , \regs[13][18] , \regs[13][17] , \regs[13][16] ,
         \regs[13][15] , \regs[13][14] , \regs[13][13] , \regs[13][12] ,
         \regs[13][11] , \regs[13][10] , \regs[13][9] , \regs[13][8] ,
         \regs[13][7] , \regs[13][6] , \regs[13][5] , \regs[13][4] ,
         \regs[13][3] , \regs[13][2] , \regs[13][1] , \regs[13][0] ,
         \regs[14][31] , \regs[14][30] , \regs[14][29] , \regs[14][28] ,
         \regs[14][27] , \regs[14][26] , \regs[14][25] , \regs[14][24] ,
         \regs[14][23] , \regs[14][22] , \regs[14][21] , \regs[14][20] ,
         \regs[14][19] , \regs[14][18] , \regs[14][17] , \regs[14][16] ,
         \regs[14][15] , \regs[14][14] , \regs[14][13] , \regs[14][12] ,
         \regs[14][11] , \regs[14][10] , \regs[14][9] , \regs[14][8] ,
         \regs[14][7] , \regs[14][6] , \regs[14][5] , \regs[14][4] ,
         \regs[14][3] , \regs[14][2] , \regs[14][1] , \regs[14][0] ,
         \regs[15][31] , \regs[15][30] , \regs[15][29] , \regs[15][28] ,
         \regs[15][27] , \regs[15][26] , \regs[15][25] , \regs[15][24] ,
         \regs[15][23] , \regs[15][22] , \regs[15][21] , \regs[15][20] ,
         \regs[15][19] , \regs[15][18] , \regs[15][17] , \regs[15][16] ,
         \regs[15][15] , \regs[15][14] , \regs[15][13] , \regs[15][12] ,
         \regs[15][11] , \regs[15][10] , \regs[15][9] , \regs[15][8] ,
         \regs[15][7] , \regs[15][6] , \regs[15][5] , \regs[15][4] ,
         \regs[15][3] , \regs[15][2] , \regs[15][1] , \regs[15][0] ,
         \regs[16][31] , \regs[16][30] , \regs[16][29] , \regs[16][28] ,
         \regs[16][27] , \regs[16][26] , \regs[16][25] , \regs[16][24] ,
         \regs[16][23] , \regs[16][22] , \regs[16][21] , \regs[16][20] ,
         \regs[16][19] , \regs[16][18] , \regs[16][17] , \regs[16][16] ,
         \regs[16][15] , \regs[16][14] , \regs[16][13] , \regs[16][12] ,
         \regs[16][11] , \regs[16][10] , \regs[16][9] , \regs[16][8] ,
         \regs[16][7] , \regs[16][6] , \regs[16][5] , \regs[16][4] ,
         \regs[16][3] , \regs[16][2] , \regs[16][1] , \regs[16][0] ,
         \regs[17][31] , \regs[17][30] , \regs[17][29] , \regs[17][28] ,
         \regs[17][27] , \regs[17][26] , \regs[17][25] , \regs[17][24] ,
         \regs[17][23] , \regs[17][22] , \regs[17][21] , \regs[17][20] ,
         \regs[17][19] , \regs[17][18] , \regs[17][17] , \regs[17][16] ,
         \regs[17][15] , \regs[17][14] , \regs[17][13] , \regs[17][12] ,
         \regs[17][11] , \regs[17][10] , \regs[17][9] , \regs[17][8] ,
         \regs[17][7] , \regs[17][6] , \regs[17][5] , \regs[17][4] ,
         \regs[17][3] , \regs[17][2] , \regs[17][1] , \regs[17][0] ,
         \regs[18][31] , \regs[18][30] , \regs[18][29] , \regs[18][28] ,
         \regs[18][27] , \regs[18][26] , \regs[18][25] , \regs[18][24] ,
         \regs[18][23] , \regs[18][22] , \regs[18][21] , \regs[18][20] ,
         \regs[18][19] , \regs[18][18] , \regs[18][17] , \regs[18][16] ,
         \regs[18][15] , \regs[18][14] , \regs[18][13] , \regs[18][12] ,
         \regs[18][11] , \regs[18][10] , \regs[18][9] , \regs[18][8] ,
         \regs[18][7] , \regs[18][6] , \regs[18][5] , \regs[18][4] ,
         \regs[18][3] , \regs[18][2] , \regs[18][1] , \regs[18][0] ,
         \regs[19][31] , \regs[19][30] , \regs[19][29] , \regs[19][28] ,
         \regs[19][27] , \regs[19][26] , \regs[19][25] , \regs[19][24] ,
         \regs[19][23] , \regs[19][22] , \regs[19][21] , \regs[19][20] ,
         \regs[19][19] , \regs[19][18] , \regs[19][17] , \regs[19][16] ,
         \regs[19][15] , \regs[19][14] , \regs[19][13] , \regs[19][12] ,
         \regs[19][11] , \regs[19][10] , \regs[19][9] , \regs[19][8] ,
         \regs[19][7] , \regs[19][6] , \regs[19][5] , \regs[19][4] ,
         \regs[19][3] , \regs[19][2] , \regs[19][1] , \regs[19][0] ,
         \regs[20][31] , \regs[20][30] , \regs[20][29] , \regs[20][28] ,
         \regs[20][27] , \regs[20][26] , \regs[20][25] , \regs[20][24] ,
         \regs[20][23] , \regs[20][22] , \regs[20][21] , \regs[20][20] ,
         \regs[20][19] , \regs[20][18] , \regs[20][17] , \regs[20][16] ,
         \regs[20][15] , \regs[20][14] , \regs[20][13] , \regs[20][12] ,
         \regs[20][11] , \regs[20][10] , \regs[20][9] , \regs[20][8] ,
         \regs[20][7] , \regs[20][6] , \regs[20][5] , \regs[20][4] ,
         \regs[20][3] , \regs[20][2] , \regs[20][1] , \regs[20][0] ,
         \regs[21][31] , \regs[21][30] , \regs[21][29] , \regs[21][28] ,
         \regs[21][27] , \regs[21][26] , \regs[21][25] , \regs[21][24] ,
         \regs[21][23] , \regs[21][22] , \regs[21][21] , \regs[21][20] ,
         \regs[21][19] , \regs[21][18] , \regs[21][17] , \regs[21][16] ,
         \regs[21][15] , \regs[21][14] , \regs[21][13] , \regs[21][12] ,
         \regs[21][11] , \regs[21][10] , \regs[21][9] , \regs[21][8] ,
         \regs[21][7] , \regs[21][6] , \regs[21][5] , \regs[21][4] ,
         \regs[21][3] , \regs[21][2] , \regs[21][1] , \regs[21][0] ,
         \regs[22][31] , \regs[22][30] , \regs[22][29] , \regs[22][28] ,
         \regs[22][27] , \regs[22][26] , \regs[22][25] , \regs[22][24] ,
         \regs[22][23] , \regs[22][22] , \regs[22][21] , \regs[22][20] ,
         \regs[22][19] , \regs[22][18] , \regs[22][17] , \regs[22][16] ,
         \regs[22][15] , \regs[22][14] , \regs[22][13] , \regs[22][12] ,
         \regs[22][11] , \regs[22][10] , \regs[22][9] , \regs[22][8] ,
         \regs[22][7] , \regs[22][6] , \regs[22][5] , \regs[22][4] ,
         \regs[22][3] , \regs[22][2] , \regs[22][1] , \regs[22][0] ,
         \regs[23][31] , \regs[23][30] , \regs[23][29] , \regs[23][28] ,
         \regs[23][27] , \regs[23][26] , \regs[23][25] , \regs[23][24] ,
         \regs[23][23] , \regs[23][22] , \regs[23][21] , \regs[23][20] ,
         \regs[23][19] , \regs[23][18] , \regs[23][17] , \regs[23][16] ,
         \regs[23][15] , \regs[23][14] , \regs[23][13] , \regs[23][12] ,
         \regs[23][11] , \regs[23][10] , \regs[23][9] , \regs[23][8] ,
         \regs[23][7] , \regs[23][6] , \regs[23][5] , \regs[23][4] ,
         \regs[23][3] , \regs[23][2] , \regs[23][1] , \regs[23][0] ,
         \regs[24][31] , \regs[24][30] , \regs[24][29] , \regs[24][28] ,
         \regs[24][27] , \regs[24][26] , \regs[24][25] , \regs[24][24] ,
         \regs[24][23] , \regs[24][22] , \regs[24][21] , \regs[24][20] ,
         \regs[24][19] , \regs[24][18] , \regs[24][17] , \regs[24][16] ,
         \regs[24][15] , \regs[24][14] , \regs[24][13] , \regs[24][12] ,
         \regs[24][11] , \regs[24][10] , \regs[24][9] , \regs[24][8] ,
         \regs[24][7] , \regs[24][6] , \regs[24][5] , \regs[24][4] ,
         \regs[24][3] , \regs[24][2] , \regs[24][1] , \regs[24][0] ,
         \regs[25][31] , \regs[25][30] , \regs[25][29] , \regs[25][28] ,
         \regs[25][27] , \regs[25][26] , \regs[25][25] , \regs[25][24] ,
         \regs[25][23] , \regs[25][22] , \regs[25][21] , \regs[25][20] ,
         \regs[25][19] , \regs[25][18] , \regs[25][17] , \regs[25][16] ,
         \regs[25][15] , \regs[25][14] , \regs[25][13] , \regs[25][12] ,
         \regs[25][11] , \regs[25][10] , \regs[25][9] , \regs[25][8] ,
         \regs[25][7] , \regs[25][6] , \regs[25][5] , \regs[25][4] ,
         \regs[25][3] , \regs[25][2] , \regs[25][1] , \regs[25][0] ,
         \regs[26][31] , \regs[26][30] , \regs[26][29] , \regs[26][28] ,
         \regs[26][27] , \regs[26][26] , \regs[26][25] , \regs[26][24] ,
         \regs[26][23] , \regs[26][22] , \regs[26][21] , \regs[26][20] ,
         \regs[26][19] , \regs[26][18] , \regs[26][17] , \regs[26][16] ,
         \regs[26][15] , \regs[26][14] , \regs[26][13] , \regs[26][12] ,
         \regs[26][11] , \regs[26][10] , \regs[26][9] , \regs[26][8] ,
         \regs[26][7] , \regs[26][6] , \regs[26][5] , \regs[26][4] ,
         \regs[26][3] , \regs[26][2] , \regs[26][1] , \regs[26][0] ,
         \regs[27][31] , \regs[27][30] , \regs[27][29] , \regs[27][28] ,
         \regs[27][27] , \regs[27][26] , \regs[27][25] , \regs[27][24] ,
         \regs[27][23] , \regs[27][22] , \regs[27][21] , \regs[27][20] ,
         \regs[27][19] , \regs[27][18] , \regs[27][17] , \regs[27][16] ,
         \regs[27][15] , \regs[27][14] , \regs[27][13] , \regs[27][12] ,
         \regs[27][11] , \regs[27][10] , \regs[27][9] , \regs[27][8] ,
         \regs[27][7] , \regs[27][6] , \regs[27][5] , \regs[27][4] ,
         \regs[27][3] , \regs[27][2] , \regs[27][1] , \regs[27][0] ,
         \regs[28][31] , \regs[28][30] , \regs[28][29] , \regs[28][28] ,
         \regs[28][27] , \regs[28][26] , \regs[28][25] , \regs[28][24] ,
         \regs[28][23] , \regs[28][22] , \regs[28][21] , \regs[28][20] ,
         \regs[28][19] , \regs[28][18] , \regs[28][17] , \regs[28][16] ,
         \regs[28][15] , \regs[28][14] , \regs[28][13] , \regs[28][12] ,
         \regs[28][11] , \regs[28][10] , \regs[28][9] , \regs[28][8] ,
         \regs[28][7] , \regs[28][6] , \regs[28][5] , \regs[28][4] ,
         \regs[28][3] , \regs[28][2] , \regs[28][1] , \regs[28][0] ,
         \regs[29][31] , \regs[29][30] , \regs[29][29] , \regs[29][28] ,
         \regs[29][27] , \regs[29][26] , \regs[29][25] , \regs[29][24] ,
         \regs[29][23] , \regs[29][22] , \regs[29][21] , \regs[29][20] ,
         \regs[29][19] , \regs[29][18] , \regs[29][17] , \regs[29][16] ,
         \regs[29][15] , \regs[29][14] , \regs[29][13] , \regs[29][12] ,
         \regs[29][11] , \regs[29][10] , \regs[29][9] , \regs[29][8] ,
         \regs[29][7] , \regs[29][6] , \regs[29][5] , \regs[29][4] ,
         \regs[29][3] , \regs[29][2] , \regs[29][1] , \regs[29][0] ,
         \regs[30][31] , \regs[30][30] , \regs[30][29] , \regs[30][28] ,
         \regs[30][27] , \regs[30][26] , \regs[30][25] , \regs[30][24] ,
         \regs[30][23] , \regs[30][22] , \regs[30][21] , \regs[30][20] ,
         \regs[30][19] , \regs[30][18] , \regs[30][17] , \regs[30][16] ,
         \regs[30][15] , \regs[30][14] , \regs[30][13] , \regs[30][12] ,
         \regs[30][11] , \regs[30][10] , \regs[30][9] , \regs[30][8] ,
         \regs[30][7] , \regs[30][6] , \regs[30][5] , \regs[30][4] ,
         \regs[30][3] , \regs[30][2] , \regs[30][1] , \regs[30][0] ,
         \regs[31][31] , \regs[31][30] , \regs[31][29] , \regs[31][28] ,
         \regs[31][27] , \regs[31][26] , \regs[31][25] , \regs[31][24] ,
         \regs[31][23] , \regs[31][22] , \regs[31][21] , \regs[31][20] ,
         \regs[31][19] , \regs[31][18] , \regs[31][17] , \regs[31][16] ,
         \regs[31][15] , \regs[31][14] , \regs[31][13] , \regs[31][12] ,
         \regs[31][11] , \regs[31][10] , \regs[31][9] , \regs[31][8] ,
         \regs[31][7] , \regs[31][6] , \regs[31][5] , \regs[31][4] ,
         \regs[31][3] , \regs[31][2] , \regs[31][1] , \regs[31][0] , n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n82, n84, n85, n86, n87, n88,
         n89, n90, n91, n93, n94, n95, n96, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n113, n116, n117, n118, n119,
         n120, n122, n125, n126, n127, n128, n129, n130, n131, n132, n135,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n150, n152, n153, n154, n155, n160, n161, n162, n163, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n192, n193, n194, n195, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n220, n221, n222, n223, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n336, n337, n338, n339, n340, n341,
         n342, n343, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n459, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n511, n512, n513, n514,
         n515, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n636, n637, n639, n640, n641,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n670, n671, n672, n673, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n692, n693, n694, n695, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n718, n719, n720, n721, n722, n723, n724, n725, n726, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n820, n821,
         n823, n824, n825, n827, n828, n829, n830, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n848,
         n852, n855, n857, n858, n859, n865, n866, n867, n868, n874, n875,
         n876, n877, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n894, n899, n902, n904, n905, n906, n915, n916, n917, n918,
         n927, n928, n929, n930, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n950, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n985, n986, n987, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n1000, n1001, n1002, n1003, n1004, n1005,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1040, n1042, n1043, n1044, n1045, n1048, n1049, n1050,
         n1051, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1071, n1073, n1074, n1075,
         n1076, n1081, n1082, n1083, n1084, n1089, n1090, n1091, n1092, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1112, n1114, n1115, n1116, n1117, n1123, n1124, n1125, n1126, n1130,
         n1131, n1132, n1133, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1157, n1158, n1159, n1160, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1210, n1211, n1212, n1213, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2688, n2689, n2690, n2691, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2740, n2742, n2743, n2744, n2745, n2750, n2751, n2752, n2753, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2771, n2773, n2774, n2775, n2776, n2779,
         n2780, n2781, n2782, n2787, n2788, n2789, n2790, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2809, n2811,
         n2813, n2814, n2815, n2819, n2820, n2821, n2822, n2829, n2830, n2831,
         n2832, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2852, n2855, n2857, n2858, n2859, n2868, n2869, n2870,
         n2871, n2880, n2881, n2882, n2883, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2905, n2914, n2955, n2956,
         n2965, n2974, n2983, n2992, n2993, n3002, n3003, n3012, n3021, n3030,
         n3031, n3040, n3049, n3058, n3067, n3068, n3077, n3078, n3087, n3096,
         n3105, n3106, n3115, n3124, n3133, n3142, n3143, n3154, n3163, n3172,
         n3181, n3182, n3191, n3192, n3193, n3202, n3203, n3212, n3213, n3254,
         n3255, n3256, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503;

  DFFX1_LVT \regs_reg[4][30]  ( .D(n2433), .CLK(clk), .Q(\regs[4][30] ) );
  DFFX1_LVT \regs_reg[16][31]  ( .D(n2050), .CLK(clk), .Q(\regs[16][31] ) );
  DFFX1_LVT \regs_reg[23][31]  ( .D(n1826), .CLK(clk), .Q(\regs[23][31] ) );
  DFFX1_LVT \regs_reg[30][30]  ( .D(n1601), .CLK(clk), .Q(\regs[30][30] ) );
  DFFX1_LVT \regs_reg[8][30]  ( .D(n2305), .CLK(clk), .Q(\regs[8][30] ) );
  DFFX1_LVT \regs_reg[20][31]  ( .D(n1922), .CLK(clk), .Q(\regs[20][31] ) );
  DFFX1_LVT \regs_reg[12][30]  ( .D(n2177), .CLK(clk), .Q(\regs[12][30] ) );
  DFFX1_LVT \regs_reg[16][29]  ( .D(n2048), .CLK(clk), .Q(\regs[16][29] ) );
  DFFX1_LVT \regs_reg[19][30]  ( .D(n1953), .CLK(clk), .Q(\regs[19][30] ) );
  DFFX1_LVT \regs_reg[22][29]  ( .D(n1856), .CLK(clk), .Q(\regs[22][29] ) );
  DFFX1_LVT \regs_reg[23][30]  ( .D(n1825), .CLK(clk), .Q(\regs[23][30] ) );
  DFFX1_LVT \regs_reg[16][30]  ( .D(n2049), .CLK(clk), .Q(\regs[16][30] ) );
  DFFX1_LVT \regs_reg[20][30]  ( .D(n1921), .CLK(clk), .Q(\regs[20][30] ) );
  DFFX1_LVT \regs_reg[3][30]  ( .D(n2465), .CLK(clk), .Q(\regs[3][30] ) );
  DFFX1_LVT \regs_reg[22][31]  ( .D(n1858), .CLK(clk), .Q(\regs[22][31] ) );
  DFFX1_LVT \regs_reg[19][31]  ( .D(n1954), .CLK(clk), .Q(\regs[19][31] ) );
  DFFX1_LVT \regs_reg[28][30]  ( .D(n1665), .CLK(clk), .Q(\regs[28][30] ) );
  DFFX1_LVT \regs_reg[11][30]  ( .D(n2209), .CLK(clk), .Q(\regs[11][30] ) );
  DFFX1_LVT \regs_reg[4][31]  ( .D(n2434), .CLK(clk), .Q(\regs[4][31] ) );
  DFFX1_LVT \regs_reg[30][31]  ( .D(n1602), .CLK(clk), .Q(\regs[30][31] ) );
  DFFX1_LVT \regs_reg[18][31]  ( .D(n1986), .CLK(clk), .Q(\regs[18][31] ) );
  DFFX1_LVT \regs_reg[6][31]  ( .D(n2370), .CLK(clk), .Q(\regs[6][31] ) );
  DFFX1_LVT \regs_reg[27][31]  ( .D(n1698), .CLK(clk), .Q(\regs[27][31] ) );
  DFFX1_LVT \regs_reg[11][31]  ( .D(n2210), .CLK(clk), .Q(\regs[11][31] ) );
  DFFX1_LVT \regs_reg[25][30]  ( .D(n1761), .CLK(clk), .Q(\regs[25][30] ) );
  DFFX1_LVT \regs_reg[22][30]  ( .D(n1857), .CLK(clk), .Q(\regs[22][30] ) );
  DFFX1_LVT \regs_reg[28][31]  ( .D(n1666), .CLK(clk), .Q(\regs[28][31] ) );
  DFFX1_LVT \regs_reg[10][31]  ( .D(n2242), .CLK(clk), .Q(\regs[10][31] ) );
  DFFX1_LVT \regs_reg[1][29]  ( .D(n2528), .CLK(clk), .Q(\regs[1][29] ) );
  DFFX1_LVT \regs_reg[12][31]  ( .D(n2178), .CLK(clk), .Q(\regs[12][31] ) );
  DFFX1_LVT \regs_reg[10][29]  ( .D(n2240), .CLK(clk), .Q(\regs[10][29] ) );
  DFFX1_LVT \regs_reg[11][28]  ( .D(n2207), .CLK(clk), .Q(\regs[11][28] ) );
  DFFX1_LVT \regs_reg[22][28]  ( .D(n1855), .CLK(clk), .Q(\regs[22][28] ) );
  DFFX1_LVT \regs_reg[13][29]  ( .D(n2144), .CLK(clk), .Q(\regs[13][29] ) );
  DFFX1_LVT \regs_reg[17][29]  ( .D(n2016), .CLK(clk), .Q(\regs[17][29] ) );
  DFFX1_LVT \regs_reg[14][29]  ( .D(n2112), .CLK(clk), .Q(\regs[14][29] ) );
  DFFX1_LVT \regs_reg[18][29]  ( .D(n1984), .CLK(clk), .Q(\regs[18][29] ) );
  DFFX1_LVT \regs_reg[8][29]  ( .D(n2304), .CLK(clk), .Q(\regs[8][29] ) );
  DFFX1_LVT \regs_reg[11][29]  ( .D(n2208), .CLK(clk), .Q(\regs[11][29] ) );
  DFFX1_LVT \regs_reg[20][29]  ( .D(n1920), .CLK(clk), .Q(\regs[20][29] ) );
  DFFX1_LVT \regs_reg[18][28]  ( .D(n1983), .CLK(clk), .Q(\regs[18][28] ) );
  DFFX1_LVT \regs_reg[19][29]  ( .D(n1952), .CLK(clk), .Q(\regs[19][29] ) );
  DFFX1_LVT \regs_reg[19][28]  ( .D(n1951), .CLK(clk), .Q(\regs[19][28] ) );
  DFFX1_LVT \regs_reg[28][27]  ( .D(n1662), .CLK(clk), .Q(\regs[28][27] ) );
  DFFX1_LVT \regs_reg[13][28]  ( .D(n2143), .CLK(clk), .Q(\regs[13][28] ) );
  DFFX1_LVT \regs_reg[27][28]  ( .D(n1695), .CLK(clk), .Q(\regs[27][28] ) );
  DFFX1_LVT \regs_reg[30][28]  ( .D(n1599), .CLK(clk), .Q(\regs[30][28] ) );
  DFFX1_LVT \regs_reg[25][28]  ( .D(n1759), .CLK(clk), .Q(\regs[25][28] ) );
  DFFX1_LVT \regs_reg[4][28]  ( .D(n2431), .CLK(clk), .Q(\regs[4][28] ) );
  DFFX1_LVT \regs_reg[20][28]  ( .D(n1919), .CLK(clk), .Q(\regs[20][28] ) );
  DFFX1_LVT \regs_reg[11][27]  ( .D(n2206), .CLK(clk), .Q(\regs[11][27] ) );
  DFFX1_LVT \regs_reg[25][27]  ( .D(n1758), .CLK(clk), .Q(\regs[25][27] ) );
  DFFX1_LVT \regs_reg[16][28]  ( .D(n2047), .CLK(clk), .Q(\regs[16][28] ) );
  DFFX1_LVT \regs_reg[28][28]  ( .D(n1663), .CLK(clk), .Q(\regs[28][28] ) );
  DFFX1_LVT \regs_reg[13][27]  ( .D(n2142), .CLK(clk), .Q(\regs[13][27] ) );
  DFFX1_LVT \regs_reg[20][26]  ( .D(n1917), .CLK(clk), .Q(\regs[20][26] ) );
  DFFX1_LVT \regs_reg[4][27]  ( .D(n2430), .CLK(clk), .Q(\regs[4][27] ) );
  DFFX1_LVT \regs_reg[12][27]  ( .D(n2174), .CLK(clk), .Q(\regs[12][27] ) );
  DFFX1_LVT \regs_reg[18][27]  ( .D(n1982), .CLK(clk), .Q(\regs[18][27] ) );
  DFFX1_LVT \regs_reg[1][27]  ( .D(n2526), .CLK(clk), .Q(\regs[1][27] ) );
  DFFX1_LVT \regs_reg[19][27]  ( .D(n1950), .CLK(clk), .Q(\regs[19][27] ) );
  DFFX1_LVT \regs_reg[3][27]  ( .D(n2462), .CLK(clk), .Q(\regs[3][27] ) );
  DFFX1_LVT \regs_reg[30][27]  ( .D(n1598), .CLK(clk), .Q(\regs[30][27] ) );
  DFFX1_LVT \regs_reg[7][27]  ( .D(n2334), .CLK(clk), .Q(\regs[7][27] ) );
  DFFX1_LVT \regs_reg[9][27]  ( .D(n2270), .CLK(clk), .Q(\regs[9][27] ) );
  DFFX1_LVT \regs_reg[16][27]  ( .D(n2046), .CLK(clk), .Q(\regs[16][27] ) );
  DFFX1_LVT \regs_reg[18][26]  ( .D(n1981), .CLK(clk), .Q(\regs[18][26] ) );
  DFFX1_LVT \regs_reg[22][27]  ( .D(n1854), .CLK(clk), .Q(\regs[22][27] ) );
  DFFX1_LVT \regs_reg[17][27]  ( .D(n2014), .CLK(clk), .Q(\regs[17][27] ) );
  DFFX1_LVT \regs_reg[6][27]  ( .D(n2366), .CLK(clk), .Q(\regs[6][27] ) );
  DFFX1_LVT \regs_reg[19][26]  ( .D(n1949), .CLK(clk), .Q(\regs[19][26] ) );
  DFFX1_LVT \regs_reg[7][26]  ( .D(n2333), .CLK(clk), .Q(\regs[7][26] ) );
  DFFX1_LVT \regs_reg[16][26]  ( .D(n2045), .CLK(clk), .Q(\regs[16][26] ) );
  DFFX1_LVT \regs_reg[4][26]  ( .D(n2429), .CLK(clk), .Q(\regs[4][26] ) );
  DFFX1_LVT \regs_reg[27][26]  ( .D(n1693), .CLK(clk), .Q(\regs[27][26] ) );
  DFFX1_LVT \regs_reg[28][26]  ( .D(n1661), .CLK(clk), .Q(\regs[28][26] ) );
  DFFX1_LVT \regs_reg[3][26]  ( .D(n2461), .CLK(clk), .Q(\regs[3][26] ) );
  DFFX1_LVT \regs_reg[25][26]  ( .D(n1757), .CLK(clk), .Q(\regs[25][26] ) );
  DFFX1_LVT \regs_reg[6][26]  ( .D(n2365), .CLK(clk), .Q(\regs[6][26] ) );
  DFFX1_LVT \regs_reg[22][26]  ( .D(n1853), .CLK(clk), .Q(\regs[22][26] ) );
  DFFX1_LVT \regs_reg[9][26]  ( .D(n2269), .CLK(clk), .Q(\regs[9][26] ) );
  DFFX1_LVT \regs_reg[23][26]  ( .D(n1821), .CLK(clk), .Q(\regs[23][26] ) );
  DFFX1_LVT \regs_reg[11][26]  ( .D(n2205), .CLK(clk), .Q(\regs[11][26] ) );
  DFFX1_LVT \regs_reg[16][25]  ( .D(n2044), .CLK(clk), .Q(\regs[16][25] ) );
  DFFX1_LVT \regs_reg[14][24]  ( .D(n2107), .CLK(clk), .Q(\regs[14][24] ) );
  DFFX1_LVT \regs_reg[6][25]  ( .D(n2364), .CLK(clk), .Q(\regs[6][25] ) );
  DFFX1_LVT \regs_reg[13][24]  ( .D(n2139), .CLK(clk), .Q(\regs[13][24] ) );
  DFFX1_LVT \regs_reg[20][25]  ( .D(n1916), .CLK(clk), .Q(\regs[20][25] ) );
  DFFX1_LVT \regs_reg[19][25]  ( .D(n1948), .CLK(clk), .Q(\regs[19][25] ) );
  DFFX1_LVT \regs_reg[8][25]  ( .D(n2300), .CLK(clk), .Q(\regs[8][25] ) );
  DFFX1_LVT \regs_reg[14][25]  ( .D(n2108), .CLK(clk), .Q(\regs[14][25] ) );
  DFFX1_LVT \regs_reg[11][25]  ( .D(n2204), .CLK(clk), .Q(\regs[11][25] ) );
  DFFX1_LVT \regs_reg[4][25]  ( .D(n2428), .CLK(clk), .Q(\regs[4][25] ) );
  DFFX1_LVT \regs_reg[12][25]  ( .D(n2172), .CLK(clk), .Q(\regs[12][25] ) );
  DFFX1_LVT \regs_reg[4][24]  ( .D(n2427), .CLK(clk), .Q(\regs[4][24] ) );
  DFFX1_LVT \regs_reg[23][24]  ( .D(n1819), .CLK(clk), .Q(\regs[23][24] ) );
  DFFX1_LVT \regs_reg[9][25]  ( .D(n2268), .CLK(clk), .Q(\regs[9][25] ) );
  DFFX1_LVT \regs_reg[27][25]  ( .D(n1692), .CLK(clk), .Q(\regs[27][25] ) );
  DFFX1_LVT \regs_reg[20][24]  ( .D(n1915), .CLK(clk), .Q(\regs[20][24] ) );
  DFFX1_LVT \regs_reg[3][24]  ( .D(n2459), .CLK(clk), .Q(\regs[3][24] ) );
  DFFX1_LVT \regs_reg[4][23]  ( .D(n2426), .CLK(clk), .Q(\regs[4][23] ) );
  DFFX1_LVT \regs_reg[18][24]  ( .D(n1979), .CLK(clk), .Q(\regs[18][24] ) );
  DFFX1_LVT \regs_reg[22][24]  ( .D(n1851), .CLK(clk), .Q(\regs[22][24] ) );
  DFFX1_LVT \regs_reg[19][24]  ( .D(n1947), .CLK(clk), .Q(\regs[19][24] ) );
  DFFX1_LVT \regs_reg[29][24]  ( .D(n1627), .CLK(clk), .Q(\regs[29][24] ) );
  DFFX1_LVT \regs_reg[7][24]  ( .D(n2331), .CLK(clk), .Q(\regs[7][24] ) );
  DFFX1_LVT \regs_reg[8][24]  ( .D(n2299), .CLK(clk), .Q(\regs[8][24] ) );
  DFFX1_LVT \regs_reg[24][24]  ( .D(n1787), .CLK(clk), .Q(\regs[24][24] ) );
  DFFX1_LVT \regs_reg[6][24]  ( .D(n2363), .CLK(clk), .Q(\regs[6][24] ) );
  DFFX1_LVT \regs_reg[12][24]  ( .D(n2171), .CLK(clk), .Q(\regs[12][24] ) );
  DFFX1_LVT \regs_reg[27][24]  ( .D(n1691), .CLK(clk), .Q(\regs[27][24] ) );
  DFFX1_LVT \regs_reg[11][24]  ( .D(n2203), .CLK(clk), .Q(\regs[11][24] ) );
  DFFX1_LVT \regs_reg[20][23]  ( .D(n1914), .CLK(clk), .Q(\regs[20][23] ) );
  DFFX1_LVT \regs_reg[16][24]  ( .D(n2043), .CLK(clk), .Q(\regs[16][24] ) );
  DFFX1_LVT \regs_reg[9][24]  ( .D(n2267), .CLK(clk), .Q(\regs[9][24] ) );
  DFFX1_LVT \regs_reg[10][24]  ( .D(n2235), .CLK(clk), .Q(\regs[10][24] ) );
  DFFX1_LVT \regs_reg[20][22]  ( .D(n1913), .CLK(clk), .Q(\regs[20][22] ) );
  DFFX1_LVT \regs_reg[26][23]  ( .D(n1722), .CLK(clk), .Q(\regs[26][23] ) );
  DFFX1_LVT \regs_reg[27][23]  ( .D(n1690), .CLK(clk), .Q(\regs[27][23] ) );
  DFFX1_LVT \regs_reg[29][22]  ( .D(n1625), .CLK(clk), .Q(\regs[29][22] ) );
  DFFX1_LVT \regs_reg[14][23]  ( .D(n2106), .CLK(clk), .Q(\regs[14][23] ) );
  DFFX1_LVT \regs_reg[3][23]  ( .D(n2458), .CLK(clk), .Q(\regs[3][23] ) );
  DFFX1_LVT \regs_reg[16][23]  ( .D(n2042), .CLK(clk), .Q(\regs[16][23] ) );
  DFFX1_LVT \regs_reg[24][23]  ( .D(n1786), .CLK(clk), .Q(\regs[24][23] ) );
  DFFX1_LVT \regs_reg[11][23]  ( .D(n2202), .CLK(clk), .Q(\regs[11][23] ) );
  DFFX1_LVT \regs_reg[8][23]  ( .D(n2298), .CLK(clk), .Q(\regs[8][23] ) );
  DFFX1_LVT \regs_reg[31][23]  ( .D(n1562), .CLK(clk), .Q(\regs[31][23] ) );
  DFFX1_LVT \regs_reg[12][23]  ( .D(n2170), .CLK(clk), .Q(\regs[12][23] ) );
  DFFX1_LVT \regs_reg[9][23]  ( .D(n2266), .CLK(clk), .Q(\regs[9][23] ) );
  DFFX1_LVT \regs_reg[18][23]  ( .D(n1978), .CLK(clk), .Q(\regs[18][23] ) );
  DFFX1_LVT \regs_reg[15][22]  ( .D(n2073), .CLK(clk), .Q(\regs[15][22] ) );
  DFFX1_LVT \regs_reg[22][23]  ( .D(n1850), .CLK(clk), .Q(\regs[22][23] ) );
  DFFX1_LVT \regs_reg[31][22]  ( .D(n1561), .CLK(clk), .Q(\regs[31][22] ) );
  DFFX1_LVT \regs_reg[9][21]  ( .D(n2264), .CLK(clk), .Q(\regs[9][21] ) );
  DFFX1_LVT \regs_reg[13][22]  ( .D(n2137), .CLK(clk), .Q(\regs[13][22] ) );
  DFFX1_LVT \regs_reg[19][21]  ( .D(n1944), .CLK(clk), .Q(\regs[19][21] ) );
  DFFX1_LVT \regs_reg[6][22]  ( .D(n2361), .CLK(clk), .Q(\regs[6][22] ) );
  DFFX1_LVT \regs_reg[4][21]  ( .D(n2424), .CLK(clk), .Q(\regs[4][21] ) );
  DFFX1_LVT \regs_reg[28][22]  ( .D(n1657), .CLK(clk), .Q(\regs[28][22] ) );
  DFFX1_LVT \regs_reg[7][22]  ( .D(n2329), .CLK(clk), .Q(\regs[7][22] ) );
  DFFX1_LVT \regs_reg[23][22]  ( .D(n1817), .CLK(clk), .Q(\regs[23][22] ) );
  DFFX1_LVT \regs_reg[9][22]  ( .D(n2265), .CLK(clk), .Q(\regs[9][22] ) );
  DFFX1_LVT \regs_reg[24][22]  ( .D(n1785), .CLK(clk), .Q(\regs[24][22] ) );
  DFFX1_LVT \regs_reg[4][22]  ( .D(n2425), .CLK(clk), .Q(\regs[4][22] ) );
  DFFX1_LVT \regs_reg[11][22]  ( .D(n2201), .CLK(clk), .Q(\regs[11][22] ) );
  DFFX1_LVT \regs_reg[19][22]  ( .D(n1945), .CLK(clk), .Q(\regs[19][22] ) );
  DFFX1_LVT \regs_reg[12][22]  ( .D(n2169), .CLK(clk), .Q(\regs[12][22] ) );
  DFFX1_LVT \regs_reg[8][22]  ( .D(n2297), .CLK(clk), .Q(\regs[8][22] ) );
  DFFX1_LVT \regs_reg[16][22]  ( .D(n2041), .CLK(clk), .Q(\regs[16][22] ) );
  DFFX1_LVT \regs_reg[10][22]  ( .D(n2233), .CLK(clk), .Q(\regs[10][22] ) );
  DFFX1_LVT \regs_reg[3][22]  ( .D(n2457), .CLK(clk), .Q(\regs[3][22] ) );
  DFFX1_LVT \regs_reg[8][21]  ( .D(n2296), .CLK(clk), .Q(\regs[8][21] ) );
  DFFX1_LVT \regs_reg[18][22]  ( .D(n1977), .CLK(clk), .Q(\regs[18][22] ) );
  DFFX1_LVT \regs_reg[14][22]  ( .D(n2105), .CLK(clk), .Q(\regs[14][22] ) );
  DFFX1_LVT \regs_reg[18][20]  ( .D(n1975), .CLK(clk), .Q(\regs[18][20] ) );
  DFFX1_LVT \regs_reg[1][21]  ( .D(n2520), .CLK(clk), .Q(\regs[1][21] ) );
  DFFX1_LVT \regs_reg[16][20]  ( .D(n2039), .CLK(clk), .Q(\regs[16][20] ) );
  DFFX1_LVT \regs_reg[3][21]  ( .D(n2456), .CLK(clk), .Q(\regs[3][21] ) );
  DFFX1_LVT \regs_reg[9][20]  ( .D(n2263), .CLK(clk), .Q(\regs[9][20] ) );
  DFFX1_LVT \regs_reg[21][21]  ( .D(n1880), .CLK(clk), .Q(\regs[21][21] ) );
  DFFX1_LVT \regs_reg[5][21]  ( .D(n2392), .CLK(clk), .Q(\regs[5][21] ) );
  DFFX1_LVT \regs_reg[18][21]  ( .D(n1976), .CLK(clk), .Q(\regs[18][21] ) );
  DFFX1_LVT \regs_reg[16][21]  ( .D(n2040), .CLK(clk), .Q(\regs[16][21] ) );
  DFFX1_LVT \regs_reg[30][21]  ( .D(n1592), .CLK(clk), .Q(\regs[30][21] ) );
  DFFX1_LVT \regs_reg[25][21]  ( .D(n1752), .CLK(clk), .Q(\regs[25][21] ) );
  DFFX1_LVT \regs_reg[10][21]  ( .D(n2232), .CLK(clk), .Q(\regs[10][21] ) );
  DFFX1_LVT \regs_reg[22][21]  ( .D(n1848), .CLK(clk), .Q(\regs[22][21] ) );
  DFFX1_LVT \regs_reg[12][21]  ( .D(n2168), .CLK(clk), .Q(\regs[12][21] ) );
  DFFX1_LVT \regs_reg[27][21]  ( .D(n1688), .CLK(clk), .Q(\regs[27][21] ) );
  DFFX1_LVT \regs_reg[11][20]  ( .D(n2199), .CLK(clk), .Q(\regs[11][20] ) );
  DFFX1_LVT \regs_reg[3][20]  ( .D(n2455), .CLK(clk), .Q(\regs[3][20] ) );
  DFFX1_LVT \regs_reg[15][21]  ( .D(n2072), .CLK(clk), .Q(\regs[15][21] ) );
  DFFX1_LVT \regs_reg[6][21]  ( .D(n2360), .CLK(clk), .Q(\regs[6][21] ) );
  DFFX1_LVT \regs_reg[11][21]  ( .D(n2200), .CLK(clk), .Q(\regs[11][21] ) );
  DFFX1_LVT \regs_reg[4][20]  ( .D(n2423), .CLK(clk), .Q(\regs[4][20] ) );
  DFFX1_LVT \regs_reg[8][20]  ( .D(n2295), .CLK(clk), .Q(\regs[8][20] ) );
  DFFX1_LVT \regs_reg[30][20]  ( .D(n1591), .CLK(clk), .Q(\regs[30][20] ) );
  DFFX1_LVT \regs_reg[24][20]  ( .D(n1783), .CLK(clk), .Q(\regs[24][20] ) );
  DFFX1_LVT \regs_reg[6][20]  ( .D(n2359), .CLK(clk), .Q(\regs[6][20] ) );
  DFFX1_LVT \regs_reg[28][20]  ( .D(n1655), .CLK(clk), .Q(\regs[28][20] ) );
  DFFX1_LVT \regs_reg[31][20]  ( .D(n1559), .CLK(clk), .Q(\regs[31][20] ) );
  DFFX1_LVT \regs_reg[14][20]  ( .D(n2103), .CLK(clk), .Q(\regs[14][20] ) );
  DFFX1_LVT \regs_reg[12][20]  ( .D(n2167), .CLK(clk), .Q(\regs[12][20] ) );
  DFFX1_LVT \regs_reg[25][20]  ( .D(n1751), .CLK(clk), .Q(\regs[25][20] ) );
  DFFX1_LVT \regs_reg[13][20]  ( .D(n2135), .CLK(clk), .Q(\regs[13][20] ) );
  DFFX1_LVT \regs_reg[27][20]  ( .D(n1687), .CLK(clk), .Q(\regs[27][20] ) );
  DFFX1_LVT \regs_reg[19][20]  ( .D(n1943), .CLK(clk), .Q(\regs[19][20] ) );
  DFFX1_LVT \regs_reg[20][20]  ( .D(n1911), .CLK(clk), .Q(\regs[20][20] ) );
  DFFX1_LVT \regs_reg[8][18]  ( .D(n2293), .CLK(clk), .Q(\regs[8][18] ) );
  DFFX1_LVT \regs_reg[7][18]  ( .D(n2325), .CLK(clk), .Q(\regs[7][18] ) );
  DFFX1_LVT \regs_reg[11][18]  ( .D(n2197), .CLK(clk), .Q(\regs[11][18] ) );
  DFFX1_LVT \regs_reg[6][19]  ( .D(n2358), .CLK(clk), .Q(\regs[6][19] ) );
  DFFX1_LVT \regs_reg[16][19]  ( .D(n2038), .CLK(clk), .Q(\regs[16][19] ) );
  DFFX1_LVT \regs_reg[21][19]  ( .D(n1878), .CLK(clk), .Q(\regs[21][19] ) );
  DFFX1_LVT \regs_reg[3][19]  ( .D(n2454), .CLK(clk), .Q(\regs[3][19] ) );
  DFFX1_LVT \regs_reg[13][19]  ( .D(n2134), .CLK(clk), .Q(\regs[13][19] ) );
  DFFX1_LVT \regs_reg[9][19]  ( .D(n2262), .CLK(clk), .Q(\regs[9][19] ) );
  DFFX1_LVT \regs_reg[31][19]  ( .D(n1558), .CLK(clk), .Q(\regs[31][19] ) );
  DFFX1_LVT \regs_reg[10][19]  ( .D(n2230), .CLK(clk), .Q(\regs[10][19] ) );
  DFFX1_LVT \regs_reg[14][19]  ( .D(n2102), .CLK(clk), .Q(\regs[14][19] ) );
  DFFX1_LVT \regs_reg[25][19]  ( .D(n1750), .CLK(clk), .Q(\regs[25][19] ) );
  DFFX1_LVT \regs_reg[23][19]  ( .D(n1814), .CLK(clk), .Q(\regs[23][19] ) );
  DFFX1_LVT \regs_reg[8][19]  ( .D(n2294), .CLK(clk), .Q(\regs[8][19] ) );
  DFFX1_LVT \regs_reg[18][18]  ( .D(n1973), .CLK(clk), .Q(\regs[18][18] ) );
  DFFX1_LVT \regs_reg[19][19]  ( .D(n1942), .CLK(clk), .Q(\regs[19][19] ) );
  DFFX1_LVT \regs_reg[30][19]  ( .D(n1590), .CLK(clk), .Q(\regs[30][19] ) );
  DFFX1_LVT \regs_reg[11][19]  ( .D(n2198), .CLK(clk), .Q(\regs[11][19] ) );
  DFFX1_LVT \regs_reg[24][19]  ( .D(n1782), .CLK(clk), .Q(\regs[24][19] ) );
  DFFX1_LVT \regs_reg[20][18]  ( .D(n1909), .CLK(clk), .Q(\regs[20][18] ) );
  DFFX1_LVT \regs_reg[27][17]  ( .D(n1684), .CLK(clk), .Q(\regs[27][17] ) );
  DFFX1_LVT \regs_reg[20][17]  ( .D(n1908), .CLK(clk), .Q(\regs[20][17] ) );
  DFFX1_LVT \regs_reg[9][17]  ( .D(n2260), .CLK(clk), .Q(\regs[9][17] ) );
  DFFX1_LVT \regs_reg[19][18]  ( .D(n1941), .CLK(clk), .Q(\regs[19][18] ) );
  DFFX1_LVT \regs_reg[6][18]  ( .D(n2357), .CLK(clk), .Q(\regs[6][18] ) );
  DFFX1_LVT \regs_reg[13][18]  ( .D(n2133), .CLK(clk), .Q(\regs[13][18] ) );
  DFFX1_LVT \regs_reg[3][18]  ( .D(n2453), .CLK(clk), .Q(\regs[3][18] ) );
  DFFX1_LVT \regs_reg[15][18]  ( .D(n2069), .CLK(clk), .Q(\regs[15][18] ) );
  DFFX1_LVT \regs_reg[12][18]  ( .D(n2165), .CLK(clk), .Q(\regs[12][18] ) );
  DFFX1_LVT \regs_reg[5][18]  ( .D(n2389), .CLK(clk), .Q(\regs[5][18] ) );
  DFFX1_LVT \regs_reg[21][18]  ( .D(n1877), .CLK(clk), .Q(\regs[21][18] ) );
  DFFX1_LVT \regs_reg[28][18]  ( .D(n1653), .CLK(clk), .Q(\regs[28][18] ) );
  DFFX1_LVT \regs_reg[4][18]  ( .D(n2421), .CLK(clk), .Q(\regs[4][18] ) );
  DFFX1_LVT \regs_reg[16][18]  ( .D(n2037), .CLK(clk), .Q(\regs[16][18] ) );
  DFFX1_LVT \regs_reg[3][17]  ( .D(n2452), .CLK(clk), .Q(\regs[3][17] ) );
  DFFX1_LVT \regs_reg[31][18]  ( .D(n1557), .CLK(clk), .Q(\regs[31][18] ) );
  DFFX1_LVT \regs_reg[17][18]  ( .D(n2005), .CLK(clk), .Q(\regs[17][18] ) );
  DFFX1_LVT \regs_reg[27][18]  ( .D(n1685), .CLK(clk), .Q(\regs[27][18] ) );
  DFFX1_LVT \regs_reg[14][18]  ( .D(n2101), .CLK(clk), .Q(\regs[14][18] ) );
  DFFX1_LVT \regs_reg[15][17]  ( .D(n2068), .CLK(clk), .Q(\regs[15][17] ) );
  DFFX1_LVT \regs_reg[29][16]  ( .D(n1619), .CLK(clk), .Q(\regs[29][16] ) );
  DFFX1_LVT \regs_reg[5][17]  ( .D(n2388), .CLK(clk), .Q(\regs[5][17] ) );
  DFFX1_LVT \regs_reg[19][17]  ( .D(n1940), .CLK(clk), .Q(\regs[19][17] ) );
  DFFX1_LVT \regs_reg[25][17]  ( .D(n1748), .CLK(clk), .Q(\regs[25][17] ) );
  DFFX1_LVT \regs_reg[11][17]  ( .D(n2196), .CLK(clk), .Q(\regs[11][17] ) );
  DFFX1_LVT \regs_reg[30][17]  ( .D(n1588), .CLK(clk), .Q(\regs[30][17] ) );
  DFFX1_LVT \regs_reg[10][17]  ( .D(n2228), .CLK(clk), .Q(\regs[10][17] ) );
  DFFX1_LVT \regs_reg[7][17]  ( .D(n2324), .CLK(clk), .Q(\regs[7][17] ) );
  DFFX1_LVT \regs_reg[1][17]  ( .D(n2516), .CLK(clk), .Q(\regs[1][17] ) );
  DFFX1_LVT \regs_reg[16][17]  ( .D(n2036), .CLK(clk), .Q(\regs[16][17] ) );
  DFFX1_LVT \regs_reg[12][16]  ( .D(n2163), .CLK(clk), .Q(\regs[12][16] ) );
  DFFX1_LVT \regs_reg[12][17]  ( .D(n2164), .CLK(clk), .Q(\regs[12][17] ) );
  DFFX1_LVT \regs_reg[31][17]  ( .D(n1556), .CLK(clk), .Q(\regs[31][17] ) );
  DFFX1_LVT \regs_reg[18][17]  ( .D(n1972), .CLK(clk), .Q(\regs[18][17] ) );
  DFFX1_LVT \regs_reg[13][17]  ( .D(n2132), .CLK(clk), .Q(\regs[13][17] ) );
  DFFX1_LVT \regs_reg[4][17]  ( .D(n2420), .CLK(clk), .Q(\regs[4][17] ) );
  DFFX1_LVT \regs_reg[30][15]  ( .D(n1586), .CLK(clk), .Q(\regs[30][15] ) );
  DFFX1_LVT \regs_reg[15][16]  ( .D(n2067), .CLK(clk), .Q(\regs[15][16] ) );
  DFFX1_LVT \regs_reg[20][16]  ( .D(n1907), .CLK(clk), .Q(\regs[20][16] ) );
  DFFX1_LVT \regs_reg[23][16]  ( .D(n1811), .CLK(clk), .Q(\regs[23][16] ) );
  DFFX1_LVT \regs_reg[6][16]  ( .D(n2355), .CLK(clk), .Q(\regs[6][16] ) );
  DFFX1_LVT \regs_reg[9][16]  ( .D(n2259), .CLK(clk), .Q(\regs[9][16] ) );
  DFFX1_LVT \regs_reg[8][16]  ( .D(n2291), .CLK(clk), .Q(\regs[8][16] ) );
  DFFX1_LVT \regs_reg[4][16]  ( .D(n2419), .CLK(clk), .Q(\regs[4][16] ) );
  DFFX1_LVT \regs_reg[3][16]  ( .D(n2451), .CLK(clk), .Q(\regs[3][16] ) );
  DFFX1_LVT \regs_reg[11][16]  ( .D(n2195), .CLK(clk), .Q(\regs[11][16] ) );
  DFFX1_LVT \regs_reg[14][16]  ( .D(n2099), .CLK(clk), .Q(\regs[14][16] ) );
  DFFX1_LVT \regs_reg[18][16]  ( .D(n1971), .CLK(clk), .Q(\regs[18][16] ) );
  DFFX1_LVT \regs_reg[16][15]  ( .D(n2034), .CLK(clk), .Q(\regs[16][15] ) );
  DFFX1_LVT \regs_reg[16][16]  ( .D(n2035), .CLK(clk), .Q(\regs[16][16] ) );
  DFFX1_LVT \regs_reg[22][16]  ( .D(n1843), .CLK(clk), .Q(\regs[22][16] ) );
  DFFX1_LVT \regs_reg[4][15]  ( .D(n2418), .CLK(clk), .Q(\regs[4][15] ) );
  DFFX1_LVT \regs_reg[8][15]  ( .D(n2290), .CLK(clk), .Q(\regs[8][15] ) );
  DFFX1_LVT \regs_reg[23][14]  ( .D(n1809), .CLK(clk), .Q(\regs[23][14] ) );
  DFFX1_LVT \regs_reg[3][15]  ( .D(n2450), .CLK(clk), .Q(\regs[3][15] ) );
  DFFX1_LVT \regs_reg[6][15]  ( .D(n2354), .CLK(clk), .Q(\regs[6][15] ) );
  DFFX1_LVT \regs_reg[7][15]  ( .D(n2322), .CLK(clk), .Q(\regs[7][15] ) );
  DFFX1_LVT \regs_reg[12][15]  ( .D(n2162), .CLK(clk), .Q(\regs[12][15] ) );
  DFFX1_LVT \regs_reg[25][15]  ( .D(n1746), .CLK(clk), .Q(\regs[25][15] ) );
  DFFX1_LVT \regs_reg[14][15]  ( .D(n2098), .CLK(clk), .Q(\regs[14][15] ) );
  DFFX1_LVT \regs_reg[11][15]  ( .D(n2194), .CLK(clk), .Q(\regs[11][15] ) );
  DFFX1_LVT \regs_reg[23][15]  ( .D(n1810), .CLK(clk), .Q(\regs[23][15] ) );
  DFFX1_LVT \regs_reg[28][15]  ( .D(n1650), .CLK(clk), .Q(\regs[28][15] ) );
  DFFX1_LVT \regs_reg[18][15]  ( .D(n1970), .CLK(clk), .Q(\regs[18][15] ) );
  DFFX1_LVT \regs_reg[20][15]  ( .D(n1906), .CLK(clk), .Q(\regs[20][15] ) );
  DFFX1_LVT \regs_reg[29][15]  ( .D(n1618), .CLK(clk), .Q(\regs[29][15] ) );
  DFFX1_LVT \regs_reg[4][13]  ( .D(n2416), .CLK(clk), .Q(\regs[4][13] ) );
  DFFX1_LVT \regs_reg[29][13]  ( .D(n1616), .CLK(clk), .Q(\regs[29][13] ) );
  DFFX1_LVT \regs_reg[12][14]  ( .D(n2161), .CLK(clk), .Q(\regs[12][14] ) );
  DFFX1_LVT \regs_reg[16][14]  ( .D(n2033), .CLK(clk), .Q(\regs[16][14] ) );
  DFFX1_LVT \regs_reg[7][14]  ( .D(n2321), .CLK(clk), .Q(\regs[7][14] ) );
  DFFX1_LVT \regs_reg[14][14]  ( .D(n2097), .CLK(clk), .Q(\regs[14][14] ) );
  DFFX1_LVT \regs_reg[11][14]  ( .D(n2193), .CLK(clk), .Q(\regs[11][14] ) );
  DFFX1_LVT \regs_reg[4][14]  ( .D(n2417), .CLK(clk), .Q(\regs[4][14] ) );
  DFFX1_LVT \regs_reg[9][14]  ( .D(n2257), .CLK(clk), .Q(\regs[9][14] ) );
  DFFX1_LVT \regs_reg[30][14]  ( .D(n1585), .CLK(clk), .Q(\regs[30][14] ) );
  DFFX1_LVT \regs_reg[20][14]  ( .D(n1905), .CLK(clk), .Q(\regs[20][14] ) );
  DFFX1_LVT \regs_reg[11][13]  ( .D(n2192), .CLK(clk), .Q(\regs[11][13] ) );
  DFFX1_LVT \regs_reg[1][13]  ( .D(n2512), .CLK(clk), .Q(\regs[1][13] ) );
  DFFX1_LVT \regs_reg[29][12]  ( .D(n1615), .CLK(clk), .Q(\regs[29][12] ) );
  DFFX1_LVT \regs_reg[18][13]  ( .D(n1968), .CLK(clk), .Q(\regs[18][13] ) );
  DFFX1_LVT \regs_reg[19][13]  ( .D(n1936), .CLK(clk), .Q(\regs[19][13] ) );
  DFFX1_LVT \regs_reg[7][13]  ( .D(n2320), .CLK(clk), .Q(\regs[7][13] ) );
  DFFX1_LVT \regs_reg[23][13]  ( .D(n1808), .CLK(clk), .Q(\regs[23][13] ) );
  DFFX1_LVT \regs_reg[3][13]  ( .D(n2448), .CLK(clk), .Q(\regs[3][13] ) );
  DFFX1_LVT \regs_reg[12][13]  ( .D(n2160), .CLK(clk), .Q(\regs[12][13] ) );
  DFFX1_LVT \regs_reg[13][13]  ( .D(n2128), .CLK(clk), .Q(\regs[13][13] ) );
  DFFX1_LVT \regs_reg[6][13]  ( .D(n2352), .CLK(clk), .Q(\regs[6][13] ) );
  DFFX1_LVT \regs_reg[4][12]  ( .D(n2415), .CLK(clk), .Q(\regs[4][12] ) );
  DFFX1_LVT \regs_reg[18][12]  ( .D(n1967), .CLK(clk), .Q(\regs[18][12] ) );
  DFFX1_LVT \regs_reg[14][13]  ( .D(n2096), .CLK(clk), .Q(\regs[14][13] ) );
  DFFX1_LVT \regs_reg[8][13]  ( .D(n2288), .CLK(clk), .Q(\regs[8][13] ) );
  DFFX1_LVT \regs_reg[22][13]  ( .D(n1840), .CLK(clk), .Q(\regs[22][13] ) );
  DFFX1_LVT \regs_reg[25][13]  ( .D(n1744), .CLK(clk), .Q(\regs[25][13] ) );
  DFFX1_LVT \regs_reg[16][13]  ( .D(n2032), .CLK(clk), .Q(\regs[16][13] ) );
  DFFX1_LVT \regs_reg[19][12]  ( .D(n1935), .CLK(clk), .Q(\regs[19][12] ) );
  DFFX1_LVT \regs_reg[7][11]  ( .D(n2318), .CLK(clk), .Q(\regs[7][11] ) );
  DFFX1_LVT \regs_reg[18][11]  ( .D(n1966), .CLK(clk), .Q(\regs[18][11] ) );
  DFFX1_LVT \regs_reg[22][11]  ( .D(n1838), .CLK(clk), .Q(\regs[22][11] ) );
  DFFX1_LVT \regs_reg[6][12]  ( .D(n2351), .CLK(clk), .Q(\regs[6][12] ) );
  DFFX1_LVT \regs_reg[8][12]  ( .D(n2287), .CLK(clk), .Q(\regs[8][12] ) );
  DFFX1_LVT \regs_reg[7][12]  ( .D(n2319), .CLK(clk), .Q(\regs[7][12] ) );
  DFFX1_LVT \regs_reg[30][12]  ( .D(n1583), .CLK(clk), .Q(\regs[30][12] ) );
  DFFX1_LVT \regs_reg[16][12]  ( .D(n2031), .CLK(clk), .Q(\regs[16][12] ) );
  DFFX1_LVT \regs_reg[23][12]  ( .D(n1807), .CLK(clk), .Q(\regs[23][12] ) );
  DFFX1_LVT \regs_reg[25][12]  ( .D(n1743), .CLK(clk), .Q(\regs[25][12] ) );
  DFFX1_LVT \regs_reg[10][12]  ( .D(n2223), .CLK(clk), .Q(\regs[10][12] ) );
  DFFX1_LVT \regs_reg[22][12]  ( .D(n1839), .CLK(clk), .Q(\regs[22][12] ) );
  DFFX1_LVT \regs_reg[11][12]  ( .D(n2191), .CLK(clk), .Q(\regs[11][12] ) );
  DFFX1_LVT \regs_reg[20][11]  ( .D(n1902), .CLK(clk), .Q(\regs[20][11] ) );
  DFFX1_LVT \regs_reg[14][12]  ( .D(n2095), .CLK(clk), .Q(\regs[14][12] ) );
  DFFX1_LVT \regs_reg[20][12]  ( .D(n1903), .CLK(clk), .Q(\regs[20][12] ) );
  DFFX1_LVT \regs_reg[4][11]  ( .D(n2414), .CLK(clk), .Q(\regs[4][11] ) );
  DFFX1_LVT \regs_reg[16][11]  ( .D(n2030), .CLK(clk), .Q(\regs[16][11] ) );
  DFFX1_LVT \regs_reg[23][11]  ( .D(n1806), .CLK(clk), .Q(\regs[23][11] ) );
  DFFX1_LVT \regs_reg[11][11]  ( .D(n2190), .CLK(clk), .Q(\regs[11][11] ) );
  DFFX1_LVT \regs_reg[12][11]  ( .D(n2158), .CLK(clk), .Q(\regs[12][11] ) );
  DFFX1_LVT \regs_reg[18][10]  ( .D(n1965), .CLK(clk), .Q(\regs[18][10] ) );
  DFFX1_LVT \regs_reg[11][10]  ( .D(n2189), .CLK(clk), .Q(\regs[11][10] ) );
  DFFX1_LVT \regs_reg[22][10]  ( .D(n1837), .CLK(clk), .Q(\regs[22][10] ) );
  DFFX1_LVT \regs_reg[16][10]  ( .D(n2029), .CLK(clk), .Q(\regs[16][10] ) );
  DFFX1_LVT \regs_reg[10][10]  ( .D(n2221), .CLK(clk), .Q(\regs[10][10] ) );
  DFFX1_LVT \regs_reg[30][10]  ( .D(n1581), .CLK(clk), .Q(\regs[30][10] ) );
  DFFX1_LVT \regs_reg[4][10]  ( .D(n2413), .CLK(clk), .Q(\regs[4][10] ) );
  DFFX1_LVT \regs_reg[6][10]  ( .D(n2349), .CLK(clk), .Q(\regs[6][10] ) );
  DFFX1_LVT \regs_reg[14][10]  ( .D(n2093), .CLK(clk), .Q(\regs[14][10] ) );
  DFFX1_LVT \regs_reg[9][10]  ( .D(n2253), .CLK(clk), .Q(\regs[9][10] ) );
  DFFX1_LVT \regs_reg[12][10]  ( .D(n2157), .CLK(clk), .Q(\regs[12][10] ) );
  DFFX1_LVT \regs_reg[29][10]  ( .D(n1613), .CLK(clk), .Q(\regs[29][10] ) );
  DFFX1_LVT \regs_reg[12][8]  ( .D(n2155), .CLK(clk), .Q(\regs[12][8] ) );
  DFFX1_LVT \regs_reg[20][8]  ( .D(n1899), .CLK(clk), .Q(\regs[20][8] ) );
  DFFX1_LVT \regs_reg[7][9]  ( .D(n2316), .CLK(clk), .Q(\regs[7][9] ) );
  DFFX1_LVT \regs_reg[10][9]  ( .D(n2220), .CLK(clk), .Q(\regs[10][9] ) );
  DFFX1_LVT \regs_reg[13][9]  ( .D(n2124), .CLK(clk), .Q(\regs[13][9] ) );
  DFFX1_LVT \regs_reg[14][9]  ( .D(n2092), .CLK(clk), .Q(\regs[14][9] ) );
  DFFX1_LVT \regs_reg[27][9]  ( .D(n1676), .CLK(clk), .Q(\regs[27][9] ) );
  DFFX1_LVT \regs_reg[25][9]  ( .D(n1740), .CLK(clk), .Q(\regs[25][9] ) );
  DFFX1_LVT \regs_reg[16][9]  ( .D(n2028), .CLK(clk), .Q(\regs[16][9] ) );
  DFFX1_LVT \regs_reg[6][8]  ( .D(n2347), .CLK(clk), .Q(\regs[6][8] ) );
  DFFX1_LVT \regs_reg[7][8]  ( .D(n2315), .CLK(clk), .Q(\regs[7][8] ) );
  DFFX1_LVT \regs_reg[20][9]  ( .D(n1900), .CLK(clk), .Q(\regs[20][9] ) );
  DFFX1_LVT \regs_reg[12][9]  ( .D(n2156), .CLK(clk), .Q(\regs[12][9] ) );
  DFFX1_LVT \regs_reg[28][8]  ( .D(n1643), .CLK(clk), .Q(\regs[28][8] ) );
  DFFX1_LVT \regs_reg[12][7]  ( .D(n2154), .CLK(clk), .Q(\regs[12][7] ) );
  DFFX1_LVT \regs_reg[19][7]  ( .D(n1930), .CLK(clk), .Q(\regs[19][7] ) );
  DFFX1_LVT \regs_reg[4][8]  ( .D(n2411), .CLK(clk), .Q(\regs[4][8] ) );
  DFFX1_LVT \regs_reg[16][8]  ( .D(n2027), .CLK(clk), .Q(\regs[16][8] ) );
  DFFX1_LVT \regs_reg[3][8]  ( .D(n2443), .CLK(clk), .Q(\regs[3][8] ) );
  DFFX1_LVT \regs_reg[30][8]  ( .D(n1579), .CLK(clk), .Q(\regs[30][8] ) );
  DFFX1_LVT \regs_reg[10][8]  ( .D(n2219), .CLK(clk), .Q(\regs[10][8] ) );
  DFFX1_LVT \regs_reg[11][8]  ( .D(n2187), .CLK(clk), .Q(\regs[11][8] ) );
  DFFX1_LVT \regs_reg[13][8]  ( .D(n2123), .CLK(clk), .Q(\regs[13][8] ) );
  DFFX1_LVT \regs_reg[18][8]  ( .D(n1963), .CLK(clk), .Q(\regs[18][8] ) );
  DFFX1_LVT \regs_reg[9][8]  ( .D(n2251), .CLK(clk), .Q(\regs[9][8] ) );
  DFFX1_LVT \regs_reg[3][7]  ( .D(n2442), .CLK(clk), .Q(\regs[3][7] ) );
  DFFX1_LVT \regs_reg[10][7]  ( .D(n2218), .CLK(clk), .Q(\regs[10][7] ) );
  DFFX1_LVT \regs_reg[22][8]  ( .D(n1835), .CLK(clk), .Q(\regs[22][8] ) );
  DFFX1_LVT \regs_reg[19][8]  ( .D(n1931), .CLK(clk), .Q(\regs[19][8] ) );
  DFFX1_LVT \regs_reg[31][8]  ( .D(n1547), .CLK(clk), .Q(\regs[31][8] ) );
  DFFX1_LVT \regs_reg[4][7]  ( .D(n2410), .CLK(clk), .Q(\regs[4][7] ) );
  DFFX1_LVT \regs_reg[2][7]  ( .D(n2474), .CLK(clk), .Q(\regs[2][7] ) );
  DFFX1_LVT \regs_reg[16][6]  ( .D(n2025), .CLK(clk), .Q(\regs[16][6] ) );
  DFFX1_LVT \regs_reg[15][6]  ( .D(n2057), .CLK(clk), .Q(\regs[15][6] ) );
  DFFX1_LVT \regs_reg[7][7]  ( .D(n2314), .CLK(clk), .Q(\regs[7][7] ) );
  DFFX1_LVT \regs_reg[5][7]  ( .D(n2378), .CLK(clk), .Q(\regs[5][7] ) );
  DFFX1_LVT \regs_reg[27][7]  ( .D(n1674), .CLK(clk), .Q(\regs[27][7] ) );
  DFFX1_LVT \regs_reg[13][7]  ( .D(n2122), .CLK(clk), .Q(\regs[13][7] ) );
  DFFX1_LVT \regs_reg[28][7]  ( .D(n1642), .CLK(clk), .Q(\regs[28][7] ) );
  DFFX1_LVT \regs_reg[15][7]  ( .D(n2058), .CLK(clk), .Q(\regs[15][7] ) );
  DFFX1_LVT \regs_reg[6][7]  ( .D(n2346), .CLK(clk), .Q(\regs[6][7] ) );
  DFFX1_LVT \regs_reg[18][7]  ( .D(n1962), .CLK(clk), .Q(\regs[18][7] ) );
  DFFX1_LVT \regs_reg[23][7]  ( .D(n1802), .CLK(clk), .Q(\regs[23][7] ) );
  DFFX1_LVT \regs_reg[20][7]  ( .D(n1898), .CLK(clk), .Q(\regs[20][7] ) );
  DFFX1_LVT \regs_reg[1][7]  ( .D(n2506), .CLK(clk), .Q(\regs[1][7] ) );
  DFFX1_LVT \regs_reg[4][6]  ( .D(n2409), .CLK(clk), .Q(\regs[4][6] ) );
  DFFX1_LVT \regs_reg[18][6]  ( .D(n1961), .CLK(clk), .Q(\regs[18][6] ) );
  DFFX1_LVT \regs_reg[28][6]  ( .D(n1641), .CLK(clk), .Q(\regs[28][6] ) );
  DFFX1_LVT \regs_reg[7][6]  ( .D(n2313), .CLK(clk), .Q(\regs[7][6] ) );
  DFFX1_LVT \regs_reg[20][6]  ( .D(n1897), .CLK(clk), .Q(\regs[20][6] ) );
  DFFX1_LVT \regs_reg[6][6]  ( .D(n2345), .CLK(clk), .Q(\regs[6][6] ) );
  DFFX1_LVT \regs_reg[19][6]  ( .D(n1929), .CLK(clk), .Q(\regs[19][6] ) );
  DFFX1_LVT \regs_reg[23][6]  ( .D(n1801), .CLK(clk), .Q(\regs[23][6] ) );
  DFFX1_LVT \regs_reg[12][6]  ( .D(n2153), .CLK(clk), .Q(\regs[12][6] ) );
  DFFX1_LVT \regs_reg[10][6]  ( .D(n2217), .CLK(clk), .Q(\regs[10][6] ) );
  DFFX1_LVT \regs_reg[7][5]  ( .D(n2312), .CLK(clk), .Q(\regs[7][5] ) );
  DFFX1_LVT \regs_reg[23][5]  ( .D(n1800), .CLK(clk), .Q(\regs[23][5] ) );
  DFFX1_LVT \regs_reg[15][4]  ( .D(n2055), .CLK(clk), .Q(\regs[15][4] ) );
  DFFX1_LVT \regs_reg[2][4]  ( .D(n2471), .CLK(clk), .Q(\regs[2][4] ) );
  DFFX1_LVT \regs_reg[11][5]  ( .D(n2184), .CLK(clk), .Q(\regs[11][5] ) );
  DFFX1_LVT \regs_reg[16][5]  ( .D(n2024), .CLK(clk), .Q(\regs[16][5] ) );
  DFFX1_LVT \regs_reg[20][5]  ( .D(n1896), .CLK(clk), .Q(\regs[20][5] ) );
  DFFX1_LVT \regs_reg[3][5]  ( .D(n2440), .CLK(clk), .Q(\regs[3][5] ) );
  DFFX1_LVT \regs_reg[6][5]  ( .D(n2344), .CLK(clk), .Q(\regs[6][5] ) );
  DFFX1_LVT \regs_reg[22][5]  ( .D(n1832), .CLK(clk), .Q(\regs[22][5] ) );
  DFFX1_LVT \regs_reg[27][5]  ( .D(n1672), .CLK(clk), .Q(\regs[27][5] ) );
  DFFX1_LVT \regs_reg[25][4]  ( .D(n1735), .CLK(clk), .Q(\regs[25][4] ) );
  DFFX1_LVT \regs_reg[19][5]  ( .D(n1928), .CLK(clk), .Q(\regs[19][5] ) );
  DFFX1_LVT \regs_reg[28][5]  ( .D(n1640), .CLK(clk), .Q(\regs[28][5] ) );
  DFFX1_LVT \regs_reg[12][5]  ( .D(n2152), .CLK(clk), .Q(\regs[12][5] ) );
  DFFX1_LVT \regs_reg[10][5]  ( .D(n2216), .CLK(clk), .Q(\regs[10][5] ) );
  DFFX1_LVT \regs_reg[13][4]  ( .D(n2119), .CLK(clk), .Q(\regs[13][4] ) );
  DFFX1_LVT \regs_reg[12][3]  ( .D(n2150), .CLK(clk), .Q(\regs[12][3] ) );
  DFFX1_LVT \regs_reg[11][3]  ( .D(n2182), .CLK(clk), .Q(\regs[11][3] ) );
  DFFX1_LVT \regs_reg[19][3]  ( .D(n1926), .CLK(clk), .Q(\regs[19][3] ) );
  DFFX1_LVT \regs_reg[18][4]  ( .D(n1959), .CLK(clk), .Q(\regs[18][4] ) );
  DFFX1_LVT \regs_reg[1][4]  ( .D(n2503), .CLK(clk), .Q(\regs[1][4] ) );
  DFFX1_LVT \regs_reg[27][4]  ( .D(n1671), .CLK(clk), .Q(\regs[27][4] ) );
  DFFX1_LVT \regs_reg[11][4]  ( .D(n2183), .CLK(clk), .Q(\regs[11][4] ) );
  DFFX1_LVT \regs_reg[5][4]  ( .D(n2375), .CLK(clk), .Q(\regs[5][4] ) );
  DFFX1_LVT \regs_reg[12][4]  ( .D(n2151), .CLK(clk), .Q(\regs[12][4] ) );
  DFFX1_LVT \regs_reg[17][4]  ( .D(n1991), .CLK(clk), .Q(\regs[17][4] ) );
  DFFX1_LVT \regs_reg[19][4]  ( .D(n1927), .CLK(clk), .Q(\regs[19][4] ) );
  DFFX1_LVT \regs_reg[3][4]  ( .D(n2439), .CLK(clk), .Q(\regs[3][4] ) );
  DFFX1_LVT \regs_reg[8][4]  ( .D(n2279), .CLK(clk), .Q(\regs[8][4] ) );
  DFFX1_LVT \regs_reg[6][4]  ( .D(n2343), .CLK(clk), .Q(\regs[6][4] ) );
  DFFX1_LVT \regs_reg[20][4]  ( .D(n1895), .CLK(clk), .Q(\regs[20][4] ) );
  DFFX1_LVT \regs_reg[7][4]  ( .D(n2311), .CLK(clk), .Q(\regs[7][4] ) );
  DFFX1_LVT \regs_reg[10][4]  ( .D(n2215), .CLK(clk), .Q(\regs[10][4] ) );
  DFFX1_LVT \regs_reg[22][3]  ( .D(n1830), .CLK(clk), .Q(\regs[22][3] ) );
  DFFX1_LVT \regs_reg[2][3]  ( .D(n2470), .CLK(clk), .Q(\regs[2][3] ) );
  DFFX1_LVT \regs_reg[29][2]  ( .D(n1605), .CLK(clk), .Q(\regs[29][2] ) );
  DFFX1_LVT \regs_reg[7][2]  ( .D(n2309), .CLK(clk), .Q(\regs[7][2] ) );
  DFFX1_LVT \regs_reg[8][3]  ( .D(n2278), .CLK(clk), .Q(\regs[8][3] ) );
  DFFX1_LVT \regs_reg[10][3]  ( .D(n2214), .CLK(clk), .Q(\regs[10][3] ) );
  DFFX1_LVT \regs_reg[18][3]  ( .D(n1958), .CLK(clk), .Q(\regs[18][3] ) );
  DFFX1_LVT \regs_reg[17][3]  ( .D(n1990), .CLK(clk), .Q(\regs[17][3] ) );
  DFFX1_LVT \regs_reg[9][3]  ( .D(n2246), .CLK(clk), .Q(\regs[9][3] ) );
  DFFX1_LVT \regs_reg[20][3]  ( .D(n1894), .CLK(clk), .Q(\regs[20][3] ) );
  DFFX1_LVT \regs_reg[6][3]  ( .D(n2342), .CLK(clk), .Q(\regs[6][3] ) );
  DFFX1_LVT \regs_reg[16][3]  ( .D(n2022), .CLK(clk), .Q(\regs[16][3] ) );
  DFFX1_LVT \regs_reg[28][3]  ( .D(n1638), .CLK(clk), .Q(\regs[28][3] ) );
  DFFX1_LVT \regs_reg[30][3]  ( .D(n1574), .CLK(clk), .Q(\regs[30][3] ) );
  DFFX1_LVT \regs_reg[24][3]  ( .D(n1766), .CLK(clk), .Q(\regs[24][3] ) );
  DFFX1_LVT \regs_reg[4][3]  ( .D(n2406), .CLK(clk), .Q(\regs[4][3] ) );
  DFFX1_LVT \regs_reg[31][3]  ( .D(n1542), .CLK(clk), .Q(\regs[31][3] ) );
  DFFX1_LVT \regs_reg[23][3]  ( .D(n1798), .CLK(clk), .Q(\regs[23][3] ) );
  DFFX1_LVT \regs_reg[27][3]  ( .D(n1670), .CLK(clk), .Q(\regs[27][3] ) );
  DFFX1_LVT \regs_reg[12][2]  ( .D(n2149), .CLK(clk), .Q(\regs[12][2] ) );
  DFFX1_LVT \regs_reg[21][3]  ( .D(n1862), .CLK(clk), .Q(\regs[21][3] ) );
  DFFX1_LVT \regs_reg[25][3]  ( .D(n1734), .CLK(clk), .Q(\regs[25][3] ) );
  DFFX1_LVT \regs_reg[13][3]  ( .D(n2118), .CLK(clk), .Q(\regs[13][3] ) );
  DFFX1_LVT \regs_reg[3][3]  ( .D(n2438), .CLK(clk), .Q(\regs[3][3] ) );
  DFFX1_LVT \regs_reg[15][3]  ( .D(n2054), .CLK(clk), .Q(\regs[15][3] ) );
  DFFX1_LVT \regs_reg[22][2]  ( .D(n1829), .CLK(clk), .Q(\regs[22][2] ) );
  DFFX1_LVT \regs_reg[23][2]  ( .D(n1797), .CLK(clk), .Q(\regs[23][2] ) );
  DFFX1_LVT \regs_reg[13][1]  ( .D(n2116), .CLK(clk), .Q(\regs[13][1] ) );
  DFFX1_LVT \regs_reg[14][1]  ( .D(n2084), .CLK(clk), .Q(\regs[14][1] ) );
  DFFX1_LVT \regs_reg[15][1]  ( .D(n2052), .CLK(clk), .Q(\regs[15][1] ) );
  DFFX1_LVT \regs_reg[24][2]  ( .D(n1765), .CLK(clk), .Q(\regs[24][2] ) );
  DFFX1_LVT \regs_reg[8][2]  ( .D(n2277), .CLK(clk), .Q(\regs[8][2] ) );
  DFFX1_LVT \regs_reg[19][2]  ( .D(n1925), .CLK(clk), .Q(\regs[19][2] ) );
  DFFX1_LVT \regs_reg[21][2]  ( .D(n1861), .CLK(clk), .Q(\regs[21][2] ) );
  DFFX1_LVT \regs_reg[4][2]  ( .D(n2405), .CLK(clk), .Q(\regs[4][2] ) );
  DFFX1_LVT \regs_reg[15][2]  ( .D(n2053), .CLK(clk), .Q(\regs[15][2] ) );
  DFFX1_LVT \regs_reg[6][2]  ( .D(n2341), .CLK(clk), .Q(\regs[6][2] ) );
  DFFX1_LVT \regs_reg[17][2]  ( .D(n1989), .CLK(clk), .Q(\regs[17][2] ) );
  DFFX1_LVT \regs_reg[11][2]  ( .D(n2181), .CLK(clk), .Q(\regs[11][2] ) );
  DFFX1_LVT \regs_reg[9][2]  ( .D(n2245), .CLK(clk), .Q(\regs[9][2] ) );
  DFFX1_LVT \regs_reg[25][2]  ( .D(n1733), .CLK(clk), .Q(\regs[25][2] ) );
  DFFX1_LVT \regs_reg[20][2]  ( .D(n1893), .CLK(clk), .Q(\regs[20][2] ) );
  DFFX1_LVT \regs_reg[13][2]  ( .D(n2117), .CLK(clk), .Q(\regs[13][2] ) );
  DFFX1_LVT \regs_reg[10][2]  ( .D(n2213), .CLK(clk), .Q(\regs[10][2] ) );
  DFFX1_LVT \regs_reg[28][2]  ( .D(n1637), .CLK(clk), .Q(\regs[28][2] ) );
  DFFX1_LVT \regs_reg[14][2]  ( .D(n2085), .CLK(clk), .Q(\regs[14][2] ) );
  DFFX1_LVT \regs_reg[26][2]  ( .D(n1701), .CLK(clk), .Q(\regs[26][2] ) );
  DFFX1_LVT \regs_reg[8][1]  ( .D(n2276), .CLK(clk), .Q(\regs[8][1] ) );
  DFFX1_LVT \regs_reg[22][1]  ( .D(n1828), .CLK(clk), .Q(\regs[22][1] ) );
  DFFX1_LVT \regs_reg[27][2]  ( .D(n1669), .CLK(clk), .Q(\regs[27][2] ) );
  DFFX1_LVT \regs_reg[3][2]  ( .D(n2437), .CLK(clk), .Q(\regs[3][2] ) );
  DFFX1_LVT \regs_reg[31][2]  ( .D(n1541), .CLK(clk), .Q(\regs[31][2] ) );
  DFFX1_LVT \regs_reg[9][0]  ( .D(n2243), .CLK(clk), .Q(\regs[9][0] ) );
  DFFX1_LVT \regs_reg[16][2]  ( .D(n2021), .CLK(clk), .Q(\regs[16][2] ) );
  DFFX1_LVT \regs_reg[18][2]  ( .D(n1957), .CLK(clk), .Q(\regs[18][2] ) );
  DFFX1_LVT \regs_reg[20][1]  ( .D(n1892), .CLK(clk), .Q(\regs[20][1] ) );
  DFFX1_LVT \regs_reg[1][1]  ( .D(n2500), .CLK(clk), .Q(\regs[1][1] ) );
  DFFX1_LVT \regs_reg[30][0]  ( .D(n1571), .CLK(clk), .Q(\regs[30][0] ) );
  DFFX1_LVT \regs_reg[3][0]  ( .D(n2435), .CLK(clk), .Q(\regs[3][0] ) );
  DFFX1_LVT \regs_reg[21][0]  ( .D(n1859), .CLK(clk), .Q(\regs[21][0] ) );
  DFFX1_LVT \regs_reg[29][0]  ( .D(n1603), .CLK(clk), .Q(\regs[29][0] ) );
  DFFX1_LVT \regs_reg[10][1]  ( .D(n2212), .CLK(clk), .Q(\regs[10][1] ) );
  DFFX1_LVT \regs_reg[23][1]  ( .D(n1796), .CLK(clk), .Q(\regs[23][1] ) );
  DFFX1_LVT \regs_reg[17][1]  ( .D(n1988), .CLK(clk), .Q(\regs[17][1] ) );
  DFFX1_LVT \regs_reg[7][1]  ( .D(n2308), .CLK(clk), .Q(\regs[7][1] ) );
  DFFX1_LVT \regs_reg[31][1]  ( .D(n1540), .CLK(clk), .Q(\regs[31][1] ) );
  DFFX1_LVT \regs_reg[25][1]  ( .D(n1732), .CLK(clk), .Q(\regs[25][1] ) );
  DFFX1_LVT \regs_reg[23][0]  ( .D(n1795), .CLK(clk), .Q(\regs[23][0] ) );
  DFFX1_LVT \regs_reg[10][0]  ( .D(n2211), .CLK(clk), .Q(\regs[10][0] ) );
  DFFX1_LVT \regs_reg[5][1]  ( .D(n2372), .CLK(clk), .Q(\regs[5][1] ) );
  DFFX1_LVT \regs_reg[11][1]  ( .D(n2180), .CLK(clk), .Q(\regs[11][1] ) );
  DFFX1_LVT \regs_reg[28][1]  ( .D(n1636), .CLK(clk), .Q(\regs[28][1] ) );
  DFFX1_LVT \regs_reg[18][1]  ( .D(n1956), .CLK(clk), .Q(\regs[18][1] ) );
  DFFX1_LVT \regs_reg[29][1]  ( .D(n1604), .CLK(clk), .Q(\regs[29][1] ) );
  DFFX1_LVT \regs_reg[6][1]  ( .D(n2340), .CLK(clk), .Q(\regs[6][1] ) );
  DFFX1_LVT \regs_reg[16][1]  ( .D(n2020), .CLK(clk), .Q(\regs[16][1] ) );
  DFFX1_LVT \regs_reg[12][1]  ( .D(n2148), .CLK(clk), .Q(\regs[12][1] ) );
  DFFX1_LVT \regs_reg[3][1]  ( .D(n2436), .CLK(clk), .Q(\regs[3][1] ) );
  DFFX1_LVT \regs_reg[4][1]  ( .D(n2404), .CLK(clk), .Q(\regs[4][1] ) );
  DFFX1_LVT \regs_reg[21][1]  ( .D(n1860), .CLK(clk), .Q(\regs[21][1] ) );
  DFFX1_LVT \regs_reg[26][1]  ( .D(n1700), .CLK(clk), .Q(\regs[26][1] ) );
  DFFX1_LVT \regs_reg[19][1]  ( .D(n1924), .CLK(clk), .Q(\regs[19][1] ) );
  DFFX1_LVT \regs_reg[9][1]  ( .D(n2244), .CLK(clk), .Q(\regs[9][1] ) );
  DFFX1_LVT \regs_reg[30][1]  ( .D(n1572), .CLK(clk), .Q(\regs[30][1] ) );
  DFFX1_LVT \regs_reg[2][1]  ( .D(n2468), .CLK(clk), .Q(\regs[2][1] ) );
  DFFX1_LVT \regs_reg[24][1]  ( .D(n1764), .CLK(clk), .Q(\regs[24][1] ) );
  DFFX1_LVT \regs_reg[27][1]  ( .D(n1668), .CLK(clk), .Q(\regs[27][1] ) );
  DFFX1_LVT \regs_reg[17][0]  ( .D(n1987), .CLK(clk), .Q(\regs[17][0] ) );
  DFFX1_LVT \regs_reg[24][0]  ( .D(n1763), .CLK(clk), .Q(\regs[24][0] ) );
  DFFX1_LVT \regs_reg[31][0]  ( .D(n1539), .CLK(clk), .Q(\regs[31][0] ) );
  DFFX1_LVT \regs_reg[28][0]  ( .D(n1635), .CLK(clk), .Q(\regs[28][0] ) );
  DFFX1_LVT \regs_reg[26][0]  ( .D(n1699), .CLK(clk), .Q(\regs[26][0] ) );
  DFFX1_LVT \regs_reg[11][0]  ( .D(n2179), .CLK(clk), .Q(\regs[11][0] ) );
  DFFX1_LVT \regs_reg[5][0]  ( .D(n2371), .CLK(clk), .Q(\regs[5][0] ) );
  DFFX1_LVT \regs_reg[16][0]  ( .D(n2019), .CLK(clk), .Q(\regs[16][0] ) );
  DFFX1_LVT \regs_reg[12][0]  ( .D(n2147), .CLK(clk), .Q(\regs[12][0] ) );
  DFFX1_LVT \regs_reg[13][0]  ( .D(n2115), .CLK(clk), .Q(\regs[13][0] ) );
  DFFX1_LVT \regs_reg[1][0]  ( .D(n2499), .CLK(clk), .Q(\regs[1][0] ) );
  DFFX1_LVT \regs_reg[19][0]  ( .D(n1923), .CLK(clk), .Q(\regs[19][0] ) );
  DFFX1_LVT \regs_reg[8][0]  ( .D(n2275), .CLK(clk), .Q(\regs[8][0] ) );
  DFFX1_LVT \regs_reg[22][0]  ( .D(n1827), .CLK(clk), .Q(\regs[22][0] ) );
  DFFX1_LVT \regs_reg[7][0]  ( .D(n2307), .CLK(clk), .Q(\regs[7][0] ) );
  DFFX1_LVT \regs_reg[2][0]  ( .D(n2467), .CLK(clk), .Q(\regs[2][0] ) );
  DFFX1_LVT \regs_reg[20][0]  ( .D(n1891), .CLK(clk), .Q(\regs[20][0] ) );
  DFFX1_LVT \regs_reg[6][0]  ( .D(n2339), .CLK(clk), .Q(\regs[6][0] ) );
  DFFX1_LVT \regs_reg[27][0]  ( .D(n1667), .CLK(clk), .Q(\regs[27][0] ) );
  DFFX1_LVT \regs_reg[14][0]  ( .D(n2083), .CLK(clk), .Q(\regs[14][0] ) );
  DFFX1_LVT \regs_reg[15][0]  ( .D(n2051), .CLK(clk), .Q(\regs[15][0] ) );
  DFFX1_LVT \regs_reg[25][0]  ( .D(n1731), .CLK(clk), .Q(\regs[25][0] ) );
  DFFX1_LVT \regs_reg[18][0]  ( .D(n1955), .CLK(clk), .Q(\regs[18][0] ) );
  DFFX1_LVT \regs_reg[4][0]  ( .D(n2403), .CLK(clk), .Q(\regs[4][0] ) );
  AND2X1_LVT U3 ( .A1(n3297), .A2(re2), .Y(n2) );
  INVX1_LVT U5 ( .A(raddr2[4]), .Y(n15) );
  NAND3X0_LVT U7 ( .A1(n3448), .A2(n15), .A3(n3449), .Y(n12) );
  INVX1_LVT U8 ( .A(raddr2[1]), .Y(n17) );
  INVX1_LVT U9 ( .A(raddr2[0]), .Y(n13) );
  NAND2X0_LVT U10 ( .A1(n17), .A2(n13), .Y(n10) );
  OR2X1_LVT U11 ( .A1(n12), .A2(n10), .Y(n1) );
  AND2X1_LVT U12 ( .A1(n2), .A2(n1), .Y(n77) );
  INVX1_LVT U13 ( .A(waddr[3]), .Y(n3077) );
  INVX1_LVT U14 ( .A(waddr[0]), .Y(n3191) );
  OA22X1_LVT U16 ( .A1(waddr[0]), .A2(n13), .A3(n3470), .A4(n3449), .Y(n3) );
  OA221X1_LVT U17 ( .A1(n3191), .A2(raddr2[0]), .A3(n3298), .A4(raddr2[2]), 
        .A5(n3), .Y(n6) );
  INVX1_LVT U18 ( .A(waddr[4]), .Y(n3002) );
  AO22X1_LVT U19 ( .A1(waddr[4]), .A2(raddr2[4]), .A3(n3002), .A4(n15), .Y(n5)
         );
  INVX1_LVT U20 ( .A(waddr[1]), .Y(n3192) );
  AO22X1_LVT U21 ( .A1(waddr[1]), .A2(raddr2[1]), .A3(n3192), .A4(n17), .Y(n4)
         );
  NAND4X0_LVT U22 ( .A1(we), .A2(n6), .A3(n5), .A4(n4), .Y(n7) );
  AO221X1_LVT U23 ( .A1(waddr[3]), .A2(n3448), .A3(n3077), .A4(raddr2[3]), 
        .A5(n7), .Y(n76) );
  AND3X1_LVT U27 ( .A1(raddr2[3]), .A2(raddr2[2]), .A3(n15), .Y(n41) );
  AND2X1_LVT U28 ( .A1(raddr2[1]), .A2(raddr2[0]), .Y(n57) );
  INVX1_LVT U32 ( .A(n10), .Y(n60) );
  AND3X1_LVT U33 ( .A1(raddr2[2]), .A2(n3448), .A3(n15), .Y(n27) );
  AO22X1_LVT U36 ( .A1(\regs[15][0] ), .A2(n3471), .A3(\regs[4][0] ), .A4(
        n3460), .Y(n75) );
  INVX1_LVT U40 ( .A(n12), .Y(n51) );
  AND2X1_LVT U41 ( .A1(raddr2[1]), .A2(n13), .Y(n49) );
  AO22X1_LVT U44 ( .A1(\regs[7][0] ), .A2(n3466), .A3(\regs[2][0] ), .A4(n3454), .Y(n14) );
  INVX1_LVT U45 ( .A(n14), .Y(n20) );
  AND3X1_LVT U46 ( .A1(raddr2[3]), .A2(n15), .A3(n3449), .Y(n55) );
  AND3X1_LVT U49 ( .A1(raddr2[4]), .A2(n3448), .A3(n3449), .Y(n62) );
  AO22X1_LVT U52 ( .A1(\regs[10][0] ), .A2(n3465), .A3(\regs[18][0] ), .A4(
        n3462), .Y(n16) );
  INVX1_LVT U53 ( .A(n16), .Y(n19) );
  AND2X1_LVT U54 ( .A1(raddr2[0]), .A2(n17), .Y(n64) );
  NAND2X0_LVT U57 ( .A1(\regs[5][0] ), .A2(n3455), .Y(n18) );
  NAND3X0_LVT U58 ( .A1(n20), .A2(n19), .A3(n18), .Y(n74) );
  AND3X1_LVT U62 ( .A1(raddr2[4]), .A2(raddr2[3]), .A3(n3449), .Y(n59) );
  AO22X1_LVT U66 ( .A1(\regs[30][0] ), .A2(n3473), .A3(\regs[27][0] ), .A4(
        n3484), .Y(n34) );
  AO22X1_LVT U73 ( .A1(\regs[13][0] ), .A2(n3464), .A3(\regs[14][0] ), .A4(
        n3476), .Y(n33) );
  AO22X1_LVT U80 ( .A1(\regs[19][0] ), .A2(n3456), .A3(\regs[6][0] ), .A4(
        n3479), .Y(n32) );
  AO22X1_LVT U87 ( .A1(\regs[28][0] ), .A2(n3482), .A3(\regs[25][0] ), .A4(
        n3459), .Y(n31) );
  NOR4X1_LVT U88 ( .A1(n34), .A2(n33), .A3(n32), .A4(n31), .Y(n72) );
  AND3X1_LVT U89 ( .A1(raddr2[4]), .A2(raddr2[2]), .A3(n3448), .Y(n53) );
  AO22X1_LVT U96 ( .A1(\regs[22][0] ), .A2(n3489), .A3(\regs[3][0] ), .A4(
        n3461), .Y(n48) );
  AO22X1_LVT U103 ( .A1(\regs[16][0] ), .A2(n3472), .A3(\regs[23][0] ), .A4(
        n3488), .Y(n47) );
  AO22X1_LVT U110 ( .A1(\regs[20][0] ), .A2(n3463), .A3(\regs[12][0] ), .A4(
        n3480), .Y(n46) );
  AO22X1_LVT U117 ( .A1(\regs[8][0] ), .A2(n3485), .A3(\regs[11][0] ), .A4(
        n3490), .Y(n45) );
  NOR4X1_LVT U118 ( .A1(n48), .A2(n47), .A3(n46), .A4(n45), .Y(n71) );
  AO22X1_LVT U125 ( .A1(\regs[26][0] ), .A2(n3468), .A3(\regs[1][0] ), .A4(
        n3458), .Y(n69) );
  AO22X1_LVT U132 ( .A1(\regs[21][0] ), .A2(n3477), .A3(\regs[9][0] ), .A4(
        n3457), .Y(n68) );
  AO22X1_LVT U139 ( .A1(\regs[31][0] ), .A2(n3474), .A3(\regs[24][0] ), .A4(
        n3478), .Y(n67) );
  AO22X1_LVT U146 ( .A1(\regs[17][0] ), .A2(n3467), .A3(\regs[29][0] ), .A4(
        n3487), .Y(n66) );
  NOR4X1_LVT U147 ( .A1(n69), .A2(n68), .A3(n67), .A4(n66), .Y(n70) );
  NAND3X0_LVT U148 ( .A1(n72), .A2(n71), .A3(n70), .Y(n73) );
  OR3X1_LVT U149 ( .A1(n75), .A2(n74), .A3(n73), .Y(n80) );
  INVX1_LVT U151 ( .A(n76), .Y(n78) );
  AO22X1_LVT U155 ( .A1(n8), .A2(n80), .A3(wdata[0]), .A4(n79), .Y(rdata2[0])
         );
  AO22X1_LVT U157 ( .A1(n3490), .A2(\regs[11][1] ), .A3(n3468), .A4(
        \regs[26][1] ), .Y(n108) );
  AO22X1_LVT U158 ( .A1(n3460), .A2(\regs[4][1] ), .A3(n3454), .A4(
        \regs[2][1] ), .Y(n82) );
  INVX1_LVT U159 ( .A(n82), .Y(n87) );
  AO22X1_LVT U162 ( .A1(n3476), .A2(\regs[14][1] ), .A3(n3463), .A4(
        \regs[20][1] ), .Y(n84) );
  INVX1_LVT U163 ( .A(n84), .Y(n86) );
  NAND2X0_LVT U164 ( .A1(n3484), .A2(\regs[27][1] ), .Y(n85) );
  NAND3X0_LVT U165 ( .A1(n87), .A2(n86), .A3(n85), .Y(n107) );
  AO22X1_LVT U167 ( .A1(n3488), .A2(\regs[23][1] ), .A3(n3477), .A4(
        \regs[21][1] ), .Y(n91) );
  AO22X1_LVT U168 ( .A1(n3473), .A2(\regs[30][1] ), .A3(n3459), .A4(
        \regs[25][1] ), .Y(n90) );
  AO22X1_LVT U169 ( .A1(n3471), .A2(\regs[15][1] ), .A3(n3456), .A4(
        \regs[19][1] ), .Y(n89) );
  AO22X1_LVT U171 ( .A1(n3455), .A2(\regs[5][1] ), .A3(n3474), .A4(
        \regs[31][1] ), .Y(n88) );
  NOR4X1_LVT U172 ( .A1(n91), .A2(n90), .A3(n89), .A4(n88), .Y(n105) );
  AO22X1_LVT U174 ( .A1(n3480), .A2(\regs[12][1] ), .A3(n3485), .A4(
        \regs[8][1] ), .Y(n96) );
  AO22X1_LVT U176 ( .A1(n3464), .A2(\regs[13][1] ), .A3(n3458), .A4(
        \regs[1][1] ), .Y(n95) );
  AO22X1_LVT U177 ( .A1(n3466), .A2(\regs[7][1] ), .A3(n3478), .A4(
        \regs[24][1] ), .Y(n94) );
  AO22X1_LVT U179 ( .A1(n3489), .A2(\regs[22][1] ), .A3(n3461), .A4(
        \regs[3][1] ), .Y(n93) );
  NOR4X1_LVT U180 ( .A1(n96), .A2(n95), .A3(n94), .A4(n93), .Y(n104) );
  AO22X1_LVT U182 ( .A1(n3479), .A2(\regs[6][1] ), .A3(n3457), .A4(
        \regs[9][1] ), .Y(n102) );
  AO22X1_LVT U183 ( .A1(n3462), .A2(\regs[18][1] ), .A3(n3467), .A4(
        \regs[17][1] ), .Y(n101) );
  AO22X1_LVT U185 ( .A1(n3472), .A2(\regs[16][1] ), .A3(n3487), .A4(
        \regs[29][1] ), .Y(n100) );
  AO22X1_LVT U186 ( .A1(n3465), .A2(\regs[10][1] ), .A3(n3482), .A4(
        \regs[28][1] ), .Y(n99) );
  NOR4X1_LVT U187 ( .A1(n102), .A2(n101), .A3(n100), .A4(n99), .Y(n103) );
  NAND3X0_LVT U188 ( .A1(n105), .A2(n104), .A3(n103), .Y(n106) );
  OR3X1_LVT U189 ( .A1(n108), .A2(n107), .A3(n106), .Y(n109) );
  AO22X1_LVT U191 ( .A1(n8), .A2(n109), .A3(n79), .A4(wdata[1]), .Y(rdata2[1])
         );
  AO22X1_LVT U194 ( .A1(n3462), .A2(\regs[18][2] ), .A3(n3472), .A4(
        \regs[16][2] ), .Y(n146) );
  AO22X1_LVT U196 ( .A1(n3476), .A2(\regs[14][2] ), .A3(n3489), .A4(
        \regs[22][2] ), .Y(n113) );
  INVX1_LVT U197 ( .A(n113), .Y(n119) );
  AO22X1_LVT U200 ( .A1(n3471), .A2(\regs[15][2] ), .A3(n3480), .A4(
        \regs[12][2] ), .Y(n116) );
  INVX1_LVT U201 ( .A(n116), .Y(n118) );
  NAND2X0_LVT U202 ( .A1(n3488), .A2(\regs[23][2] ), .Y(n117) );
  NAND3X0_LVT U203 ( .A1(n119), .A2(n118), .A3(n117), .Y(n145) );
  AO22X1_LVT U206 ( .A1(n3460), .A2(\regs[4][2] ), .A3(n3478), .A4(
        \regs[24][2] ), .Y(n128) );
  AO22X1_LVT U208 ( .A1(n3479), .A2(\regs[6][2] ), .A3(n3461), .A4(
        \regs[3][2] ), .Y(n127) );
  AO22X1_LVT U210 ( .A1(n3465), .A2(\regs[10][2] ), .A3(n3463), .A4(
        \regs[20][2] ), .Y(n126) );
  AO22X1_LVT U212 ( .A1(n3464), .A2(\regs[13][2] ), .A3(n3474), .A4(
        \regs[31][2] ), .Y(n125) );
  NOR4X1_LVT U213 ( .A1(n128), .A2(n127), .A3(n126), .A4(n125), .Y(n143) );
  AO22X1_LVT U215 ( .A1(n3454), .A2(\regs[2][2] ), .A3(n3457), .A4(
        \regs[9][2] ), .Y(n132) );
  AO22X1_LVT U217 ( .A1(n3482), .A2(\regs[28][2] ), .A3(n3468), .A4(
        \regs[26][2] ), .Y(n131) );
  AO22X1_LVT U220 ( .A1(n3484), .A2(\regs[27][2] ), .A3(n3458), .A4(
        \regs[1][2] ), .Y(n130) );
  AO22X1_LVT U221 ( .A1(n3459), .A2(\regs[25][2] ), .A3(n3485), .A4(
        \regs[8][2] ), .Y(n129) );
  NOR4X1_LVT U222 ( .A1(n132), .A2(n131), .A3(n130), .A4(n129), .Y(n142) );
  AO22X1_LVT U224 ( .A1(n3490), .A2(\regs[11][2] ), .A3(n3477), .A4(
        \regs[21][2] ), .Y(n140) );
  AO22X1_LVT U226 ( .A1(n3466), .A2(\regs[7][2] ), .A3(n3473), .A4(
        \regs[30][2] ), .Y(n139) );
  AO22X1_LVT U229 ( .A1(n3455), .A2(\regs[5][2] ), .A3(n3467), .A4(
        \regs[17][2] ), .Y(n138) );
  AO22X1_LVT U232 ( .A1(n3456), .A2(\regs[19][2] ), .A3(n3487), .A4(
        \regs[29][2] ), .Y(n137) );
  NOR4X1_LVT U233 ( .A1(n140), .A2(n139), .A3(n138), .A4(n137), .Y(n141) );
  NAND3X0_LVT U234 ( .A1(n143), .A2(n142), .A3(n141), .Y(n144) );
  OR3X1_LVT U235 ( .A1(n146), .A2(n145), .A3(n144), .Y(n147) );
  AO22X1_LVT U237 ( .A1(n8), .A2(n147), .A3(n79), .A4(wdata[2]), .Y(rdata2[2])
         );
  AO22X1_LVT U239 ( .A1(n3454), .A2(\regs[2][3] ), .A3(n3476), .A4(
        \regs[14][3] ), .Y(n178) );
  AO22X1_LVT U241 ( .A1(n3456), .A2(\regs[19][3] ), .A3(n3487), .A4(
        \regs[29][3] ), .Y(n150) );
  INVX1_LVT U242 ( .A(n150), .Y(n155) );
  AO22X1_LVT U244 ( .A1(n3471), .A2(\regs[15][3] ), .A3(n3488), .A4(
        \regs[23][3] ), .Y(n152) );
  INVX1_LVT U245 ( .A(n152), .Y(n154) );
  NAND2X0_LVT U246 ( .A1(n3489), .A2(\regs[22][3] ), .Y(n153) );
  NAND3X0_LVT U247 ( .A1(n155), .A2(n154), .A3(n153), .Y(n177) );
  AO22X1_LVT U249 ( .A1(n3466), .A2(\regs[7][3] ), .A3(n3461), .A4(
        \regs[3][3] ), .Y(n163) );
  AO22X1_LVT U251 ( .A1(n3477), .A2(\regs[21][3] ), .A3(n3474), .A4(
        \regs[31][3] ), .Y(n162) );
  AO22X1_LVT U252 ( .A1(n3472), .A2(\regs[16][3] ), .A3(n3467), .A4(
        \regs[17][3] ), .Y(n161) );
  AO22X1_LVT U254 ( .A1(n3482), .A2(\regs[28][3] ), .A3(n3459), .A4(
        \regs[25][3] ), .Y(n160) );
  NOR4X1_LVT U255 ( .A1(n163), .A2(n162), .A3(n161), .A4(n160), .Y(n175) );
  AO22X1_LVT U256 ( .A1(n3484), .A2(\regs[27][3] ), .A3(n3480), .A4(
        \regs[12][3] ), .Y(n168) );
  AO22X1_LVT U257 ( .A1(n3462), .A2(\regs[18][3] ), .A3(n3478), .A4(
        \regs[24][3] ), .Y(n167) );
  AO22X1_LVT U259 ( .A1(n3463), .A2(\regs[20][3] ), .A3(n3458), .A4(
        \regs[1][3] ), .Y(n166) );
  AO22X1_LVT U260 ( .A1(n3464), .A2(\regs[13][3] ), .A3(n3468), .A4(
        \regs[26][3] ), .Y(n165) );
  NOR4X1_LVT U261 ( .A1(n168), .A2(n167), .A3(n166), .A4(n165), .Y(n174) );
  AO22X1_LVT U262 ( .A1(n3460), .A2(\regs[4][3] ), .A3(n3457), .A4(
        \regs[9][3] ), .Y(n172) );
  AO22X1_LVT U263 ( .A1(n3455), .A2(\regs[5][3] ), .A3(n3473), .A4(
        \regs[30][3] ), .Y(n171) );
  AO22X1_LVT U264 ( .A1(n3465), .A2(\regs[10][3] ), .A3(n3490), .A4(
        \regs[11][3] ), .Y(n170) );
  AO22X1_LVT U265 ( .A1(n3479), .A2(\regs[6][3] ), .A3(n3485), .A4(
        \regs[8][3] ), .Y(n169) );
  NOR4X1_LVT U266 ( .A1(n172), .A2(n171), .A3(n170), .A4(n169), .Y(n173) );
  NAND3X0_LVT U267 ( .A1(n175), .A2(n174), .A3(n173), .Y(n176) );
  OR3X1_LVT U268 ( .A1(n178), .A2(n177), .A3(n176), .Y(n179) );
  AO22X1_LVT U270 ( .A1(n8), .A2(n179), .A3(n79), .A4(wdata[3]), .Y(rdata2[3])
         );
  AO22X1_LVT U271 ( .A1(n3471), .A2(\regs[15][4] ), .A3(n3468), .A4(
        \regs[26][4] ), .Y(n207) );
  AO22X1_LVT U272 ( .A1(n3465), .A2(\regs[10][4] ), .A3(n3464), .A4(
        \regs[13][4] ), .Y(n180) );
  INVX1_LVT U273 ( .A(n180), .Y(n184) );
  AO22X1_LVT U274 ( .A1(n3466), .A2(\regs[7][4] ), .A3(n3489), .A4(
        \regs[22][4] ), .Y(n181) );
  INVX1_LVT U275 ( .A(n181), .Y(n183) );
  NAND2X0_LVT U276 ( .A1(n3490), .A2(\regs[11][4] ), .Y(n182) );
  NAND3X0_LVT U277 ( .A1(n184), .A2(n183), .A3(n182), .Y(n206) );
  AO22X1_LVT U278 ( .A1(n3456), .A2(\regs[19][4] ), .A3(n3463), .A4(
        \regs[20][4] ), .Y(n188) );
  AO22X1_LVT U279 ( .A1(n3458), .A2(\regs[1][4] ), .A3(n3477), .A4(
        \regs[21][4] ), .Y(n187) );
  AO22X1_LVT U280 ( .A1(n3455), .A2(\regs[5][4] ), .A3(n3479), .A4(
        \regs[6][4] ), .Y(n186) );
  AO22X1_LVT U281 ( .A1(n3460), .A2(\regs[4][4] ), .A3(n3454), .A4(
        \regs[2][4] ), .Y(n185) );
  NOR4X1_LVT U282 ( .A1(n188), .A2(n187), .A3(n186), .A4(n185), .Y(n204) );
  AO22X1_LVT U285 ( .A1(n3459), .A2(\regs[25][4] ), .A3(n3485), .A4(
        \regs[8][4] ), .Y(n195) );
  AO22X1_LVT U287 ( .A1(n3488), .A2(\regs[23][4] ), .A3(n3474), .A4(
        \regs[31][4] ), .Y(n194) );
  AO22X1_LVT U288 ( .A1(n3482), .A2(\regs[28][4] ), .A3(n3461), .A4(
        \regs[3][4] ), .Y(n193) );
  AO22X1_LVT U289 ( .A1(n3472), .A2(\regs[16][4] ), .A3(n3467), .A4(
        \regs[17][4] ), .Y(n192) );
  NOR4X1_LVT U290 ( .A1(n195), .A2(n194), .A3(n193), .A4(n192), .Y(n203) );
  AO22X1_LVT U292 ( .A1(n3473), .A2(\regs[30][4] ), .A3(n3484), .A4(
        \regs[27][4] ), .Y(n201) );
  AO22X1_LVT U293 ( .A1(n3462), .A2(\regs[18][4] ), .A3(n3476), .A4(
        \regs[14][4] ), .Y(n200) );
  AO22X1_LVT U294 ( .A1(n3480), .A2(\regs[12][4] ), .A3(n3487), .A4(
        \regs[29][4] ), .Y(n199) );
  AO22X1_LVT U296 ( .A1(n3457), .A2(\regs[9][4] ), .A3(n3478), .A4(
        \regs[24][4] ), .Y(n198) );
  NOR4X1_LVT U297 ( .A1(n201), .A2(n200), .A3(n199), .A4(n198), .Y(n202) );
  NAND3X0_LVT U298 ( .A1(n204), .A2(n203), .A3(n202), .Y(n205) );
  OR3X1_LVT U299 ( .A1(n207), .A2(n206), .A3(n205), .Y(n208) );
  AO22X1_LVT U301 ( .A1(n8), .A2(n208), .A3(n79), .A4(wdata[4]), .Y(rdata2[4])
         );
  AO22X1_LVT U302 ( .A1(n3465), .A2(\regs[10][5] ), .A3(n3488), .A4(
        \regs[23][5] ), .Y(n234) );
  AO22X1_LVT U304 ( .A1(n3459), .A2(\regs[25][5] ), .A3(n3463), .A4(
        \regs[20][5] ), .Y(n210) );
  INVX1_LVT U305 ( .A(n210), .Y(n214) );
  AO22X1_LVT U306 ( .A1(n3455), .A2(\regs[5][5] ), .A3(n3457), .A4(
        \regs[9][5] ), .Y(n211) );
  INVX1_LVT U307 ( .A(n211), .Y(n213) );
  NAND2X0_LVT U308 ( .A1(n3484), .A2(\regs[27][5] ), .Y(n212) );
  NAND3X0_LVT U309 ( .A1(n214), .A2(n213), .A3(n212), .Y(n233) );
  AO22X1_LVT U310 ( .A1(n3471), .A2(\regs[15][5] ), .A3(n3466), .A4(
        \regs[7][5] ), .Y(n218) );
  AO22X1_LVT U311 ( .A1(n3456), .A2(\regs[19][5] ), .A3(n3482), .A4(
        \regs[28][5] ), .Y(n217) );
  AO22X1_LVT U312 ( .A1(n3468), .A2(\regs[26][5] ), .A3(n3474), .A4(
        \regs[31][5] ), .Y(n216) );
  AO22X1_LVT U313 ( .A1(n3460), .A2(\regs[4][5] ), .A3(n3464), .A4(
        \regs[13][5] ), .Y(n215) );
  NOR4X1_LVT U314 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .Y(n231) );
  AO22X1_LVT U316 ( .A1(n3473), .A2(\regs[30][5] ), .A3(n3461), .A4(
        \regs[3][5] ), .Y(n223) );
  AO22X1_LVT U317 ( .A1(n3462), .A2(\regs[18][5] ), .A3(n3487), .A4(
        \regs[29][5] ), .Y(n222) );
  AO22X1_LVT U318 ( .A1(n3479), .A2(\regs[6][5] ), .A3(n3485), .A4(
        \regs[8][5] ), .Y(n221) );
  AO22X1_LVT U319 ( .A1(n3489), .A2(\regs[22][5] ), .A3(n3480), .A4(
        \regs[12][5] ), .Y(n220) );
  NOR4X1_LVT U320 ( .A1(n223), .A2(n222), .A3(n221), .A4(n220), .Y(n230) );
  AO22X1_LVT U321 ( .A1(n3476), .A2(\regs[14][5] ), .A3(n3490), .A4(
        \regs[11][5] ), .Y(n228) );
  AO22X1_LVT U322 ( .A1(n3472), .A2(\regs[16][5] ), .A3(n3458), .A4(
        \regs[1][5] ), .Y(n227) );
  AO22X1_LVT U323 ( .A1(n3454), .A2(\regs[2][5] ), .A3(n3478), .A4(
        \regs[24][5] ), .Y(n226) );
  AO22X1_LVT U324 ( .A1(n3477), .A2(\regs[21][5] ), .A3(n3467), .A4(
        \regs[17][5] ), .Y(n225) );
  NOR4X1_LVT U325 ( .A1(n228), .A2(n227), .A3(n226), .A4(n225), .Y(n229) );
  NAND3X0_LVT U326 ( .A1(n231), .A2(n230), .A3(n229), .Y(n232) );
  OR3X1_LVT U327 ( .A1(n234), .A2(n233), .A3(n232), .Y(n235) );
  AO22X1_LVT U329 ( .A1(n8), .A2(n235), .A3(n79), .A4(wdata[5]), .Y(rdata2[5])
         );
  AO22X1_LVT U330 ( .A1(n3471), .A2(\regs[15][6] ), .A3(n3454), .A4(
        \regs[2][6] ), .Y(n259) );
  AO22X1_LVT U331 ( .A1(n3465), .A2(\regs[10][6] ), .A3(n3480), .A4(
        \regs[12][6] ), .Y(n236) );
  INVX1_LVT U332 ( .A(n236), .Y(n240) );
  AO22X1_LVT U333 ( .A1(n3456), .A2(\regs[19][6] ), .A3(n3485), .A4(
        \regs[8][6] ), .Y(n237) );
  INVX1_LVT U334 ( .A(n237), .Y(n239) );
  NAND2X0_LVT U335 ( .A1(n3466), .A2(\regs[7][6] ), .Y(n238) );
  NAND3X0_LVT U336 ( .A1(n240), .A2(n239), .A3(n238), .Y(n258) );
  AO22X1_LVT U337 ( .A1(n3455), .A2(\regs[5][6] ), .A3(n3457), .A4(
        \regs[9][6] ), .Y(n245) );
  AO22X1_LVT U338 ( .A1(n3488), .A2(\regs[23][6] ), .A3(n3487), .A4(
        \regs[29][6] ), .Y(n244) );
  AO22X1_LVT U339 ( .A1(n3460), .A2(\regs[4][6] ), .A3(n3490), .A4(
        \regs[11][6] ), .Y(n243) );
  AO22X1_LVT U340 ( .A1(n3463), .A2(\regs[20][6] ), .A3(n3467), .A4(
        \regs[17][6] ), .Y(n242) );
  NOR4X1_LVT U341 ( .A1(n245), .A2(n244), .A3(n243), .A4(n242), .Y(n256) );
  AO22X1_LVT U342 ( .A1(n3473), .A2(\regs[30][6] ), .A3(n3476), .A4(
        \regs[14][6] ), .Y(n249) );
  AO22X1_LVT U343 ( .A1(n3479), .A2(\regs[6][6] ), .A3(n3489), .A4(
        \regs[22][6] ), .Y(n248) );
  AO22X1_LVT U344 ( .A1(n3462), .A2(\regs[18][6] ), .A3(n3468), .A4(
        \regs[26][6] ), .Y(n247) );
  AO22X1_LVT U345 ( .A1(n3464), .A2(\regs[13][6] ), .A3(n3482), .A4(
        \regs[28][6] ), .Y(n246) );
  NOR4X1_LVT U346 ( .A1(n249), .A2(n248), .A3(n247), .A4(n246), .Y(n255) );
  AO22X1_LVT U347 ( .A1(n3459), .A2(\regs[25][6] ), .A3(n3461), .A4(
        \regs[3][6] ), .Y(n253) );
  AO22X1_LVT U348 ( .A1(n3458), .A2(\regs[1][6] ), .A3(n3477), .A4(
        \regs[21][6] ), .Y(n252) );
  AO22X1_LVT U349 ( .A1(n3472), .A2(\regs[16][6] ), .A3(n3478), .A4(
        \regs[24][6] ), .Y(n251) );
  AO22X1_LVT U350 ( .A1(n3484), .A2(\regs[27][6] ), .A3(n3474), .A4(
        \regs[31][6] ), .Y(n250) );
  NOR4X1_LVT U351 ( .A1(n253), .A2(n252), .A3(n251), .A4(n250), .Y(n254) );
  NAND3X0_LVT U352 ( .A1(n256), .A2(n255), .A3(n254), .Y(n257) );
  OR3X1_LVT U353 ( .A1(n259), .A2(n258), .A3(n257), .Y(n260) );
  AO22X1_LVT U355 ( .A1(n8), .A2(n260), .A3(n79), .A4(wdata[6]), .Y(rdata2[6])
         );
  AO22X1_LVT U356 ( .A1(n3463), .A2(\regs[20][7] ), .A3(n3490), .A4(
        \regs[11][7] ), .Y(n283) );
  AO22X1_LVT U357 ( .A1(n3466), .A2(\regs[7][7] ), .A3(n3476), .A4(
        \regs[14][7] ), .Y(n261) );
  INVX1_LVT U358 ( .A(n261), .Y(n265) );
  AO22X1_LVT U359 ( .A1(n3468), .A2(\regs[26][7] ), .A3(n3487), .A4(
        \regs[29][7] ), .Y(n262) );
  INVX1_LVT U360 ( .A(n262), .Y(n264) );
  NAND2X0_LVT U361 ( .A1(n3454), .A2(\regs[2][7] ), .Y(n263) );
  NAND3X0_LVT U362 ( .A1(n265), .A2(n264), .A3(n263), .Y(n282) );
  AO22X1_LVT U363 ( .A1(n3460), .A2(\regs[4][7] ), .A3(n3472), .A4(
        \regs[16][7] ), .Y(n269) );
  AO22X1_LVT U364 ( .A1(n3464), .A2(\regs[13][7] ), .A3(n3459), .A4(
        \regs[25][7] ), .Y(n268) );
  AO22X1_LVT U365 ( .A1(n3462), .A2(\regs[18][7] ), .A3(n3457), .A4(
        \regs[9][7] ), .Y(n267) );
  AO22X1_LVT U366 ( .A1(n3465), .A2(\regs[10][7] ), .A3(n3456), .A4(
        \regs[19][7] ), .Y(n266) );
  NOR4X1_LVT U367 ( .A1(n269), .A2(n268), .A3(n267), .A4(n266), .Y(n280) );
  AO22X1_LVT U368 ( .A1(n3479), .A2(\regs[6][7] ), .A3(n3482), .A4(
        \regs[28][7] ), .Y(n273) );
  AO22X1_LVT U369 ( .A1(n3458), .A2(\regs[1][7] ), .A3(n3478), .A4(
        \regs[24][7] ), .Y(n272) );
  AO22X1_LVT U370 ( .A1(n3473), .A2(\regs[30][7] ), .A3(n3484), .A4(
        \regs[27][7] ), .Y(n271) );
  AO22X1_LVT U371 ( .A1(n3471), .A2(\regs[15][7] ), .A3(n3467), .A4(
        \regs[17][7] ), .Y(n270) );
  NOR4X1_LVT U372 ( .A1(n273), .A2(n272), .A3(n271), .A4(n270), .Y(n279) );
  AO22X1_LVT U373 ( .A1(n3455), .A2(\regs[5][7] ), .A3(n3474), .A4(
        \regs[31][7] ), .Y(n277) );
  AO22X1_LVT U374 ( .A1(n3488), .A2(\regs[23][7] ), .A3(n3477), .A4(
        \regs[21][7] ), .Y(n276) );
  AO22X1_LVT U376 ( .A1(n3461), .A2(\regs[3][7] ), .A3(n3485), .A4(
        \regs[8][7] ), .Y(n275) );
  AO22X1_LVT U377 ( .A1(n3489), .A2(\regs[22][7] ), .A3(n3480), .A4(
        \regs[12][7] ), .Y(n274) );
  NOR4X1_LVT U378 ( .A1(n277), .A2(n276), .A3(n275), .A4(n274), .Y(n278) );
  NAND3X0_LVT U379 ( .A1(n280), .A2(n279), .A3(n278), .Y(n281) );
  OR3X1_LVT U380 ( .A1(n283), .A2(n282), .A3(n281), .Y(n284) );
  AO22X1_LVT U382 ( .A1(n8), .A2(n284), .A3(n79), .A4(wdata[7]), .Y(rdata2[7])
         );
  AO22X1_LVT U383 ( .A1(n3482), .A2(\regs[28][8] ), .A3(n3490), .A4(
        \regs[11][8] ), .Y(n308) );
  AO22X1_LVT U384 ( .A1(n3462), .A2(\regs[18][8] ), .A3(n3484), .A4(
        \regs[27][8] ), .Y(n285) );
  INVX1_LVT U385 ( .A(n285), .Y(n289) );
  AO22X1_LVT U386 ( .A1(n3465), .A2(\regs[10][8] ), .A3(n3454), .A4(
        \regs[2][8] ), .Y(n286) );
  INVX1_LVT U387 ( .A(n286), .Y(n288) );
  NAND2X0_LVT U388 ( .A1(n3456), .A2(\regs[19][8] ), .Y(n287) );
  NAND3X0_LVT U389 ( .A1(n289), .A2(n288), .A3(n287), .Y(n307) );
  AO22X1_LVT U390 ( .A1(n3459), .A2(\regs[25][8] ), .A3(n3480), .A4(
        \regs[12][8] ), .Y(n293) );
  AO22X1_LVT U391 ( .A1(n3471), .A2(\regs[15][8] ), .A3(n3485), .A4(
        \regs[8][8] ), .Y(n292) );
  AO22X1_LVT U392 ( .A1(n3488), .A2(\regs[23][8] ), .A3(n3487), .A4(
        \regs[29][8] ), .Y(n291) );
  AO22X1_LVT U393 ( .A1(n3466), .A2(\regs[7][8] ), .A3(n3489), .A4(
        \regs[22][8] ), .Y(n290) );
  NOR4X1_LVT U394 ( .A1(n293), .A2(n292), .A3(n291), .A4(n290), .Y(n305) );
  AO22X1_LVT U396 ( .A1(n3474), .A2(\regs[31][8] ), .A3(n3478), .A4(
        \regs[24][8] ), .Y(n298) );
  AO22X1_LVT U397 ( .A1(n3473), .A2(\regs[30][8] ), .A3(n3479), .A4(
        \regs[6][8] ), .Y(n297) );
  AO22X1_LVT U398 ( .A1(n3463), .A2(\regs[20][8] ), .A3(n3477), .A4(
        \regs[21][8] ), .Y(n296) );
  AO22X1_LVT U400 ( .A1(n3464), .A2(\regs[13][8] ), .A3(n3468), .A4(
        \regs[26][8] ), .Y(n295) );
  NOR4X1_LVT U401 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .Y(n304) );
  AO22X1_LVT U402 ( .A1(n3455), .A2(\regs[5][8] ), .A3(n3458), .A4(
        \regs[1][8] ), .Y(n302) );
  AO22X1_LVT U403 ( .A1(n3460), .A2(\regs[4][8] ), .A3(n3457), .A4(
        \regs[9][8] ), .Y(n301) );
  AO22X1_LVT U404 ( .A1(n3476), .A2(\regs[14][8] ), .A3(n3472), .A4(
        \regs[16][8] ), .Y(n300) );
  AO22X1_LVT U405 ( .A1(n3461), .A2(\regs[3][8] ), .A3(n3467), .A4(
        \regs[17][8] ), .Y(n299) );
  NOR4X1_LVT U406 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .Y(n303) );
  NAND3X0_LVT U407 ( .A1(n305), .A2(n304), .A3(n303), .Y(n306) );
  OR3X1_LVT U408 ( .A1(n308), .A2(n307), .A3(n306), .Y(n309) );
  AO22X1_LVT U410 ( .A1(n8), .A2(n309), .A3(n79), .A4(wdata[8]), .Y(rdata2[8])
         );
  AO22X1_LVT U411 ( .A1(n29), .A2(\regs[28][9] ), .A3(n3480), .A4(
        \regs[12][9] ), .Y(n332) );
  AO22X1_LVT U412 ( .A1(n3455), .A2(\regs[5][9] ), .A3(n110), .A4(
        \regs[18][9] ), .Y(n310) );
  INVX1_LVT U413 ( .A(n310), .Y(n314) );
  AO22X1_LVT U414 ( .A1(n9), .A2(\regs[15][9] ), .A3(n40), .A4(\regs[20][9] ), 
        .Y(n311) );
  INVX1_LVT U415 ( .A(n311), .Y(n313) );
  NAND2X0_LVT U416 ( .A1(n50), .A2(\regs[26][9] ), .Y(n312) );
  NAND3X0_LVT U417 ( .A1(n314), .A2(n313), .A3(n312), .Y(n331) );
  AO22X1_LVT U418 ( .A1(n23), .A2(\regs[27][9] ), .A3(n44), .A4(\regs[11][9] ), 
        .Y(n318) );
  AO22X1_LVT U419 ( .A1(n148), .A2(\regs[2][9] ), .A3(n65), .A4(\regs[29][9] ), 
        .Y(n317) );
  AO22X1_LVT U420 ( .A1(n37), .A2(\regs[3][9] ), .A3(n56), .A4(\regs[9][9] ), 
        .Y(n316) );
  AO22X1_LVT U421 ( .A1(n28), .A2(\regs[6][9] ), .A3(n54), .A4(\regs[21][9] ), 
        .Y(n315) );
  NOR4X1_LVT U422 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .Y(n329) );
  AO22X1_LVT U423 ( .A1(n3459), .A2(\regs[25][9] ), .A3(n36), .A4(
        \regs[22][9] ), .Y(n322) );
  AO22X1_LVT U424 ( .A1(n3456), .A2(\regs[19][9] ), .A3(n3488), .A4(
        \regs[23][9] ), .Y(n321) );
  AO22X1_LVT U425 ( .A1(n120), .A2(\regs[4][9] ), .A3(n63), .A4(\regs[17][9] ), 
        .Y(n320) );
  AO22X1_LVT U426 ( .A1(n122), .A2(\regs[10][9] ), .A3(n58), .A4(\regs[31][9] ), .Y(n319) );
  NOR4X1_LVT U427 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .Y(n328) );
  AO22X1_LVT U428 ( .A1(n24), .A2(\regs[13][9] ), .A3(n43), .A4(\regs[8][9] ), 
        .Y(n326) );
  AO22X1_LVT U429 ( .A1(n25), .A2(\regs[14][9] ), .A3(n38), .A4(\regs[16][9] ), 
        .Y(n325) );
  AO22X1_LVT U430 ( .A1(n11), .A2(\regs[7][9] ), .A3(n21), .A4(\regs[30][9] ), 
        .Y(n324) );
  AO22X1_LVT U431 ( .A1(n52), .A2(\regs[1][9] ), .A3(n3478), .A4(\regs[24][9] ), .Y(n323) );
  NOR4X1_LVT U432 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .Y(n327) );
  NAND3X0_LVT U433 ( .A1(n329), .A2(n328), .A3(n327), .Y(n330) );
  OR3X1_LVT U434 ( .A1(n332), .A2(n331), .A3(n330), .Y(n333) );
  AO22X1_LVT U436 ( .A1(n8), .A2(n333), .A3(n79), .A4(wdata[9]), .Y(rdata2[9])
         );
  AO22X1_LVT U437 ( .A1(n37), .A2(\regs[3][10] ), .A3(n61), .A4(\regs[24][10] ), .Y(n358) );
  AO22X1_LVT U438 ( .A1(n28), .A2(\regs[6][10] ), .A3(n54), .A4(\regs[21][10] ), .Y(n334) );
  INVX1_LVT U439 ( .A(n334), .Y(n339) );
  AO22X1_LVT U441 ( .A1(n43), .A2(\regs[8][10] ), .A3(n56), .A4(\regs[9][10] ), 
        .Y(n336) );
  INVX1_LVT U442 ( .A(n336), .Y(n338) );
  NAND2X0_LVT U443 ( .A1(n135), .A2(\regs[5][10] ), .Y(n337) );
  NAND3X0_LVT U444 ( .A1(n339), .A2(n338), .A3(n337), .Y(n357) );
  AO22X1_LVT U445 ( .A1(n3466), .A2(\regs[7][10] ), .A3(n52), .A4(
        \regs[1][10] ), .Y(n343) );
  AO22X1_LVT U446 ( .A1(n42), .A2(\regs[12][10] ), .A3(n58), .A4(
        \regs[31][10] ), .Y(n342) );
  AO22X1_LVT U447 ( .A1(n25), .A2(\regs[14][10] ), .A3(n26), .A4(
        \regs[19][10] ), .Y(n341) );
  AO22X1_LVT U448 ( .A1(n122), .A2(\regs[10][10] ), .A3(n63), .A4(
        \regs[17][10] ), .Y(n340) );
  NOR4X1_LVT U449 ( .A1(n343), .A2(n342), .A3(n341), .A4(n340), .Y(n355) );
  AO22X1_LVT U450 ( .A1(n29), .A2(\regs[28][10] ), .A3(n65), .A4(
        \regs[29][10] ), .Y(n348) );
  AO22X1_LVT U451 ( .A1(n40), .A2(\regs[20][10] ), .A3(n50), .A4(
        \regs[26][10] ), .Y(n347) );
  AO22X1_LVT U453 ( .A1(n9), .A2(\regs[15][10] ), .A3(n36), .A4(\regs[22][10] ), .Y(n346) );
  AO22X1_LVT U454 ( .A1(n21), .A2(\regs[30][10] ), .A3(n44), .A4(
        \regs[11][10] ), .Y(n345) );
  NOR4X1_LVT U455 ( .A1(n348), .A2(n347), .A3(n346), .A4(n345), .Y(n354) );
  AO22X1_LVT U456 ( .A1(n120), .A2(\regs[4][10] ), .A3(n23), .A4(
        \regs[27][10] ), .Y(n352) );
  AO22X1_LVT U457 ( .A1(n24), .A2(\regs[13][10] ), .A3(n30), .A4(
        \regs[25][10] ), .Y(n351) );
  AO22X1_LVT U458 ( .A1(n110), .A2(\regs[18][10] ), .A3(n39), .A4(
        \regs[23][10] ), .Y(n350) );
  AO22X1_LVT U459 ( .A1(n148), .A2(\regs[2][10] ), .A3(n38), .A4(
        \regs[16][10] ), .Y(n349) );
  NOR4X1_LVT U460 ( .A1(n352), .A2(n351), .A3(n350), .A4(n349), .Y(n353) );
  NAND3X0_LVT U461 ( .A1(n355), .A2(n354), .A3(n353), .Y(n356) );
  OR3X1_LVT U462 ( .A1(n358), .A2(n357), .A3(n356), .Y(n359) );
  AO22X1_LVT U464 ( .A1(n8), .A2(n359), .A3(n79), .A4(n3499), .Y(rdata2[10])
         );
  AO22X1_LVT U465 ( .A1(n148), .A2(\regs[2][11] ), .A3(n3461), .A4(
        \regs[3][11] ), .Y(n383) );
  AO22X1_LVT U466 ( .A1(n122), .A2(\regs[10][11] ), .A3(n23), .A4(
        \regs[27][11] ), .Y(n360) );
  INVX1_LVT U467 ( .A(n360), .Y(n364) );
  AO22X1_LVT U468 ( .A1(n43), .A2(\regs[8][11] ), .A3(n50), .A4(\regs[26][11] ), .Y(n361) );
  INVX1_LVT U469 ( .A(n361), .Y(n363) );
  NAND2X0_LVT U470 ( .A1(n30), .A2(\regs[25][11] ), .Y(n362) );
  NAND3X0_LVT U471 ( .A1(n364), .A2(n363), .A3(n362), .Y(n382) );
  AO22X1_LVT U472 ( .A1(n3464), .A2(\regs[13][11] ), .A3(n36), .A4(
        \regs[22][11] ), .Y(n368) );
  AO22X1_LVT U473 ( .A1(n28), .A2(\regs[6][11] ), .A3(n39), .A4(\regs[23][11] ), .Y(n367) );
  AO22X1_LVT U474 ( .A1(n21), .A2(\regs[30][11] ), .A3(n42), .A4(
        \regs[12][11] ), .Y(n366) );
  AO22X1_LVT U475 ( .A1(n3455), .A2(\regs[5][11] ), .A3(n29), .A4(
        \regs[28][11] ), .Y(n365) );
  NOR4X1_LVT U476 ( .A1(n368), .A2(n367), .A3(n366), .A4(n365), .Y(n380) );
  AO22X1_LVT U477 ( .A1(n54), .A2(\regs[21][11] ), .A3(n61), .A4(
        \regs[24][11] ), .Y(n373) );
  AO22X1_LVT U478 ( .A1(n9), .A2(\regs[15][11] ), .A3(n26), .A4(\regs[19][11] ), .Y(n372) );
  AO22X1_LVT U479 ( .A1(n38), .A2(\regs[16][11] ), .A3(n40), .A4(
        \regs[20][11] ), .Y(n371) );
  AO22X1_LVT U480 ( .A1(n58), .A2(\regs[31][11] ), .A3(n65), .A4(
        \regs[29][11] ), .Y(n370) );
  NOR4X1_LVT U481 ( .A1(n373), .A2(n372), .A3(n371), .A4(n370), .Y(n379) );
  AO22X1_LVT U482 ( .A1(n11), .A2(\regs[7][11] ), .A3(n63), .A4(\regs[17][11] ), .Y(n377) );
  AO22X1_LVT U483 ( .A1(n120), .A2(\regs[4][11] ), .A3(n56), .A4(\regs[9][11] ), .Y(n376) );
  AO22X1_LVT U484 ( .A1(n25), .A2(\regs[14][11] ), .A3(n44), .A4(
        \regs[11][11] ), .Y(n375) );
  AO22X1_LVT U485 ( .A1(n110), .A2(\regs[18][11] ), .A3(n52), .A4(
        \regs[1][11] ), .Y(n374) );
  NOR4X1_LVT U486 ( .A1(n377), .A2(n376), .A3(n375), .A4(n374), .Y(n378) );
  NAND3X0_LVT U487 ( .A1(n380), .A2(n379), .A3(n378), .Y(n381) );
  OR3X1_LVT U488 ( .A1(n383), .A2(n382), .A3(n381), .Y(n384) );
  AO22X1_LVT U490 ( .A1(n8), .A2(n384), .A3(n79), .A4(wdata[11]), .Y(
        rdata2[11]) );
  AO22X1_LVT U491 ( .A1(n30), .A2(\regs[25][12] ), .A3(n37), .A4(\regs[3][12] ), .Y(n408) );
  AO22X1_LVT U492 ( .A1(n58), .A2(\regs[31][12] ), .A3(n65), .A4(
        \regs[29][12] ), .Y(n385) );
  INVX1_LVT U493 ( .A(n385), .Y(n389) );
  AO22X1_LVT U494 ( .A1(n42), .A2(\regs[12][12] ), .A3(n61), .A4(
        \regs[24][12] ), .Y(n386) );
  INVX1_LVT U495 ( .A(n386), .Y(n388) );
  NAND2X0_LVT U496 ( .A1(n9), .A2(\regs[15][12] ), .Y(n387) );
  NAND3X0_LVT U497 ( .A1(n389), .A2(n388), .A3(n387), .Y(n407) );
  AO22X1_LVT U498 ( .A1(n148), .A2(\regs[2][12] ), .A3(n36), .A4(
        \regs[22][12] ), .Y(n394) );
  AO22X1_LVT U500 ( .A1(n25), .A2(\regs[14][12] ), .A3(n54), .A4(
        \regs[21][12] ), .Y(n393) );
  AO22X1_LVT U501 ( .A1(n21), .A2(\regs[30][12] ), .A3(n38), .A4(
        \regs[16][12] ), .Y(n392) );
  AO22X1_LVT U502 ( .A1(n26), .A2(\regs[19][12] ), .A3(n56), .A4(\regs[9][12] ), .Y(n391) );
  NOR4X1_LVT U503 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .Y(n405) );
  AO22X1_LVT U504 ( .A1(n3465), .A2(\regs[10][12] ), .A3(n52), .A4(
        \regs[1][12] ), .Y(n398) );
  AO22X1_LVT U505 ( .A1(n11), .A2(\regs[7][12] ), .A3(n28), .A4(\regs[6][12] ), 
        .Y(n397) );
  AO22X1_LVT U506 ( .A1(n3490), .A2(\regs[11][12] ), .A3(n63), .A4(
        \regs[17][12] ), .Y(n396) );
  AO22X1_LVT U507 ( .A1(n29), .A2(\regs[28][12] ), .A3(n3463), .A4(
        \regs[20][12] ), .Y(n395) );
  NOR4X1_LVT U508 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .Y(n404) );
  AO22X1_LVT U509 ( .A1(n39), .A2(\regs[23][12] ), .A3(n3485), .A4(
        \regs[8][12] ), .Y(n402) );
  AO22X1_LVT U510 ( .A1(n135), .A2(\regs[5][12] ), .A3(n120), .A4(
        \regs[4][12] ), .Y(n401) );
  AO22X1_LVT U511 ( .A1(n110), .A2(\regs[18][12] ), .A3(n23), .A4(
        \regs[27][12] ), .Y(n400) );
  AO22X1_LVT U512 ( .A1(n24), .A2(\regs[13][12] ), .A3(n50), .A4(
        \regs[26][12] ), .Y(n399) );
  NOR4X1_LVT U513 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .Y(n403) );
  NAND3X0_LVT U514 ( .A1(n405), .A2(n404), .A3(n403), .Y(n406) );
  OR3X1_LVT U515 ( .A1(n408), .A2(n407), .A3(n406), .Y(n409) );
  AO22X1_LVT U517 ( .A1(n8), .A2(n409), .A3(n79), .A4(wdata[12]), .Y(
        rdata2[12]) );
  AO22X1_LVT U518 ( .A1(n3454), .A2(\regs[2][13] ), .A3(n3489), .A4(
        \regs[22][13] ), .Y(n433) );
  AO22X1_LVT U519 ( .A1(n3484), .A2(\regs[27][13] ), .A3(n39), .A4(
        \regs[23][13] ), .Y(n410) );
  INVX1_LVT U520 ( .A(n410), .Y(n415) );
  AO22X1_LVT U521 ( .A1(n3472), .A2(\regs[16][13] ), .A3(n42), .A4(
        \regs[12][13] ), .Y(n411) );
  INVX1_LVT U522 ( .A(n411), .Y(n414) );
  NAND2X0_LVT U524 ( .A1(n3487), .A2(\regs[29][13] ), .Y(n413) );
  NAND3X0_LVT U525 ( .A1(n415), .A2(n414), .A3(n413), .Y(n432) );
  AO22X1_LVT U526 ( .A1(n3465), .A2(\regs[10][13] ), .A3(n25), .A4(
        \regs[14][13] ), .Y(n419) );
  AO22X1_LVT U527 ( .A1(n26), .A2(\regs[19][13] ), .A3(n28), .A4(\regs[6][13] ), .Y(n418) );
  AO22X1_LVT U528 ( .A1(n52), .A2(\regs[1][13] ), .A3(n63), .A4(\regs[17][13] ), .Y(n417) );
  AO22X1_LVT U529 ( .A1(n30), .A2(\regs[25][13] ), .A3(n61), .A4(
        \regs[24][13] ), .Y(n416) );
  NOR4X1_LVT U530 ( .A1(n419), .A2(n418), .A3(n417), .A4(n416), .Y(n430) );
  AO22X1_LVT U531 ( .A1(n11), .A2(\regs[7][13] ), .A3(n43), .A4(\regs[8][13] ), 
        .Y(n423) );
  AO22X1_LVT U532 ( .A1(n120), .A2(\regs[4][13] ), .A3(n110), .A4(
        \regs[18][13] ), .Y(n422) );
  AO22X1_LVT U533 ( .A1(n135), .A2(\regs[5][13] ), .A3(n9), .A4(\regs[15][13] ), .Y(n421) );
  AO22X1_LVT U534 ( .A1(n29), .A2(\regs[28][13] ), .A3(n3457), .A4(
        \regs[9][13] ), .Y(n420) );
  NOR4X1_LVT U535 ( .A1(n423), .A2(n422), .A3(n421), .A4(n420), .Y(n429) );
  AO22X1_LVT U536 ( .A1(n21), .A2(\regs[30][13] ), .A3(n24), .A4(
        \regs[13][13] ), .Y(n427) );
  AO22X1_LVT U537 ( .A1(n40), .A2(\regs[20][13] ), .A3(n54), .A4(
        \regs[21][13] ), .Y(n426) );
  AO22X1_LVT U538 ( .A1(n37), .A2(\regs[3][13] ), .A3(n50), .A4(\regs[26][13] ), .Y(n425) );
  AO22X1_LVT U539 ( .A1(n44), .A2(\regs[11][13] ), .A3(n58), .A4(
        \regs[31][13] ), .Y(n424) );
  NOR4X1_LVT U540 ( .A1(n427), .A2(n426), .A3(n425), .A4(n424), .Y(n428) );
  NAND3X0_LVT U541 ( .A1(n430), .A2(n429), .A3(n428), .Y(n431) );
  OR3X1_LVT U542 ( .A1(n433), .A2(n432), .A3(n431), .Y(n434) );
  AO22X1_LVT U544 ( .A1(n8), .A2(n434), .A3(n79), .A4(n3502), .Y(rdata2[13])
         );
  AO22X1_LVT U545 ( .A1(n30), .A2(\regs[25][14] ), .A3(n58), .A4(
        \regs[31][14] ), .Y(n457) );
  AO22X1_LVT U546 ( .A1(n39), .A2(\regs[23][14] ), .A3(n63), .A4(
        \regs[17][14] ), .Y(n435) );
  INVX1_LVT U547 ( .A(n435), .Y(n439) );
  AO22X1_LVT U548 ( .A1(n37), .A2(\regs[3][14] ), .A3(n61), .A4(\regs[24][14] ), .Y(n436) );
  INVX1_LVT U549 ( .A(n436), .Y(n438) );
  NAND2X0_LVT U550 ( .A1(n28), .A2(\regs[6][14] ), .Y(n437) );
  NAND3X0_LVT U551 ( .A1(n439), .A2(n438), .A3(n437), .Y(n456) );
  AO22X1_LVT U552 ( .A1(n3476), .A2(\regs[14][14] ), .A3(n29), .A4(
        \regs[28][14] ), .Y(n443) );
  AO22X1_LVT U553 ( .A1(n43), .A2(\regs[8][14] ), .A3(n65), .A4(\regs[29][14] ), .Y(n442) );
  AO22X1_LVT U554 ( .A1(n110), .A2(\regs[18][14] ), .A3(n23), .A4(
        \regs[27][14] ), .Y(n441) );
  AO22X1_LVT U555 ( .A1(n9), .A2(\regs[15][14] ), .A3(n38), .A4(\regs[16][14] ), .Y(n440) );
  NOR4X1_LVT U556 ( .A1(n443), .A2(n442), .A3(n441), .A4(n440), .Y(n454) );
  AO22X1_LVT U557 ( .A1(n135), .A2(\regs[5][14] ), .A3(n54), .A4(
        \regs[21][14] ), .Y(n447) );
  AO22X1_LVT U558 ( .A1(n11), .A2(\regs[7][14] ), .A3(n36), .A4(\regs[22][14] ), .Y(n446) );
  AO22X1_LVT U559 ( .A1(n40), .A2(\regs[20][14] ), .A3(n52), .A4(\regs[1][14] ), .Y(n445) );
  AO22X1_LVT U560 ( .A1(n120), .A2(\regs[4][14] ), .A3(n24), .A4(
        \regs[13][14] ), .Y(n444) );
  NOR4X1_LVT U561 ( .A1(n447), .A2(n446), .A3(n445), .A4(n444), .Y(n453) );
  AO22X1_LVT U562 ( .A1(n3473), .A2(\regs[30][14] ), .A3(n26), .A4(
        \regs[19][14] ), .Y(n451) );
  AO22X1_LVT U563 ( .A1(n148), .A2(\regs[2][14] ), .A3(n44), .A4(
        \regs[11][14] ), .Y(n450) );
  AO22X1_LVT U564 ( .A1(n50), .A2(\regs[26][14] ), .A3(n56), .A4(\regs[9][14] ), .Y(n449) );
  AO22X1_LVT U565 ( .A1(n122), .A2(\regs[10][14] ), .A3(n42), .A4(
        \regs[12][14] ), .Y(n448) );
  NOR4X1_LVT U566 ( .A1(n451), .A2(n450), .A3(n449), .A4(n448), .Y(n452) );
  NAND3X0_LVT U567 ( .A1(n454), .A2(n453), .A3(n452), .Y(n455) );
  OR3X1_LVT U568 ( .A1(n457), .A2(n456), .A3(n455), .Y(n459) );
  AO22X1_LVT U570 ( .A1(n8), .A2(n459), .A3(n79), .A4(n3498), .Y(rdata2[14])
         );
  AO22X1_LVT U572 ( .A1(n3462), .A2(\regs[18][15] ), .A3(n3482), .A4(
        \regs[28][15] ), .Y(n483) );
  AO22X1_LVT U573 ( .A1(n3473), .A2(\regs[30][15] ), .A3(n3467), .A4(
        \regs[17][15] ), .Y(n461) );
  INVX1_LVT U574 ( .A(n461), .Y(n465) );
  AO22X1_LVT U575 ( .A1(n3463), .A2(\regs[20][15] ), .A3(n3487), .A4(
        \regs[29][15] ), .Y(n462) );
  INVX1_LVT U576 ( .A(n462), .Y(n464) );
  NAND2X0_LVT U577 ( .A1(n3468), .A2(\regs[26][15] ), .Y(n463) );
  NAND3X0_LVT U578 ( .A1(n465), .A2(n464), .A3(n463), .Y(n482) );
  AO22X1_LVT U579 ( .A1(n54), .A2(\regs[21][15] ), .A3(n58), .A4(
        \regs[31][15] ), .Y(n469) );
  AO22X1_LVT U580 ( .A1(n120), .A2(\regs[4][15] ), .A3(n30), .A4(
        \regs[25][15] ), .Y(n468) );
  AO22X1_LVT U581 ( .A1(n3471), .A2(\regs[15][15] ), .A3(n148), .A4(
        \regs[2][15] ), .Y(n467) );
  AO22X1_LVT U582 ( .A1(n39), .A2(\regs[23][15] ), .A3(n56), .A4(\regs[9][15] ), .Y(n466) );
  NOR4X1_LVT U583 ( .A1(n469), .A2(n468), .A3(n467), .A4(n466), .Y(n480) );
  AO22X1_LVT U584 ( .A1(n122), .A2(\regs[10][15] ), .A3(n43), .A4(
        \regs[8][15] ), .Y(n473) );
  AO22X1_LVT U585 ( .A1(n52), .A2(\regs[1][15] ), .A3(n61), .A4(\regs[24][15] ), .Y(n472) );
  AO22X1_LVT U586 ( .A1(n28), .A2(\regs[6][15] ), .A3(n38), .A4(\regs[16][15] ), .Y(n471) );
  AO22X1_LVT U587 ( .A1(n135), .A2(\regs[5][15] ), .A3(n23), .A4(
        \regs[27][15] ), .Y(n470) );
  NOR4X1_LVT U588 ( .A1(n473), .A2(n472), .A3(n471), .A4(n470), .Y(n479) );
  AO22X1_LVT U589 ( .A1(n26), .A2(\regs[19][15] ), .A3(n3461), .A4(
        \regs[3][15] ), .Y(n477) );
  AO22X1_LVT U590 ( .A1(n24), .A2(\regs[13][15] ), .A3(n44), .A4(
        \regs[11][15] ), .Y(n476) );
  AO22X1_LVT U591 ( .A1(n25), .A2(\regs[14][15] ), .A3(n36), .A4(
        \regs[22][15] ), .Y(n475) );
  AO22X1_LVT U592 ( .A1(n11), .A2(\regs[7][15] ), .A3(n42), .A4(\regs[12][15] ), .Y(n474) );
  NOR4X1_LVT U593 ( .A1(n477), .A2(n476), .A3(n475), .A4(n474), .Y(n478) );
  NAND3X0_LVT U594 ( .A1(n480), .A2(n479), .A3(n478), .Y(n481) );
  OR3X1_LVT U595 ( .A1(n483), .A2(n482), .A3(n481), .Y(n484) );
  AO22X1_LVT U598 ( .A1(n8), .A2(n484), .A3(n79), .A4(n3495), .Y(rdata2[15])
         );
  AO22X1_LVT U599 ( .A1(n110), .A2(\regs[18][16] ), .A3(n63), .A4(
        \regs[17][16] ), .Y(n508) );
  AO22X1_LVT U600 ( .A1(n25), .A2(\regs[14][16] ), .A3(n44), .A4(
        \regs[11][16] ), .Y(n486) );
  INVX1_LVT U601 ( .A(n486), .Y(n490) );
  AO22X1_LVT U602 ( .A1(n38), .A2(\regs[16][16] ), .A3(n56), .A4(\regs[9][16] ), .Y(n487) );
  INVX1_LVT U603 ( .A(n487), .Y(n489) );
  NAND2X0_LVT U604 ( .A1(n65), .A2(\regs[29][16] ), .Y(n488) );
  NAND3X0_LVT U605 ( .A1(n490), .A2(n489), .A3(n488), .Y(n507) );
  AO22X1_LVT U606 ( .A1(n52), .A2(\regs[1][16] ), .A3(n61), .A4(\regs[24][16] ), .Y(n494) );
  AO22X1_LVT U607 ( .A1(n42), .A2(\regs[12][16] ), .A3(n43), .A4(\regs[8][16] ), .Y(n493) );
  AO22X1_LVT U608 ( .A1(n26), .A2(\regs[19][16] ), .A3(n50), .A4(
        \regs[26][16] ), .Y(n492) );
  AO22X1_LVT U609 ( .A1(n21), .A2(\regs[30][16] ), .A3(n30), .A4(
        \regs[25][16] ), .Y(n491) );
  NOR4X1_LVT U610 ( .A1(n494), .A2(n493), .A3(n492), .A4(n491), .Y(n505) );
  AO22X1_LVT U611 ( .A1(n29), .A2(\regs[28][16] ), .A3(n3474), .A4(
        \regs[31][16] ), .Y(n498) );
  AO22X1_LVT U612 ( .A1(n122), .A2(\regs[10][16] ), .A3(n24), .A4(
        \regs[13][16] ), .Y(n497) );
  AO22X1_LVT U613 ( .A1(n148), .A2(\regs[2][16] ), .A3(n3484), .A4(
        \regs[27][16] ), .Y(n496) );
  AO22X1_LVT U614 ( .A1(n37), .A2(\regs[3][16] ), .A3(n40), .A4(\regs[20][16] ), .Y(n495) );
  NOR4X1_LVT U615 ( .A1(n498), .A2(n497), .A3(n496), .A4(n495), .Y(n504) );
  AO22X1_LVT U616 ( .A1(n11), .A2(\regs[7][16] ), .A3(n39), .A4(\regs[23][16] ), .Y(n502) );
  AO22X1_LVT U617 ( .A1(n135), .A2(\regs[5][16] ), .A3(n28), .A4(\regs[6][16] ), .Y(n501) );
  AO22X1_LVT U618 ( .A1(n36), .A2(\regs[22][16] ), .A3(n3477), .A4(
        \regs[21][16] ), .Y(n500) );
  AO22X1_LVT U619 ( .A1(n9), .A2(\regs[15][16] ), .A3(n120), .A4(\regs[4][16] ), .Y(n499) );
  NOR4X1_LVT U620 ( .A1(n502), .A2(n501), .A3(n500), .A4(n499), .Y(n503) );
  NAND3X0_LVT U621 ( .A1(n505), .A2(n504), .A3(n503), .Y(n506) );
  OR3X1_LVT U622 ( .A1(n508), .A2(n507), .A3(n506), .Y(n509) );
  AO22X1_LVT U624 ( .A1(n8), .A2(n509), .A3(n79), .A4(wdata[16]), .Y(
        rdata2[16]) );
  AO22X1_LVT U626 ( .A1(n3471), .A2(\regs[15][17] ), .A3(n3467), .A4(
        \regs[17][17] ), .Y(n534) );
  AO22X1_LVT U627 ( .A1(n3464), .A2(\regs[13][17] ), .A3(n3479), .A4(
        \regs[6][17] ), .Y(n511) );
  INVX1_LVT U628 ( .A(n511), .Y(n515) );
  AO22X1_LVT U629 ( .A1(n3473), .A2(\regs[30][17] ), .A3(n3480), .A4(
        \regs[12][17] ), .Y(n512) );
  INVX1_LVT U630 ( .A(n512), .Y(n514) );
  NAND2X0_LVT U631 ( .A1(n3460), .A2(\regs[4][17] ), .Y(n513) );
  NAND3X0_LVT U632 ( .A1(n515), .A2(n514), .A3(n513), .Y(n533) );
  AO22X1_LVT U633 ( .A1(n3457), .A2(\regs[9][17] ), .A3(n3487), .A4(
        \regs[29][17] ), .Y(n520) );
  AO22X1_LVT U634 ( .A1(n3463), .A2(\regs[20][17] ), .A3(n3474), .A4(
        \regs[31][17] ), .Y(n519) );
  AO22X1_LVT U635 ( .A1(n3466), .A2(\regs[7][17] ), .A3(n3461), .A4(
        \regs[3][17] ), .Y(n518) );
  AO22X1_LVT U636 ( .A1(n3488), .A2(\regs[23][17] ), .A3(n3478), .A4(
        \regs[24][17] ), .Y(n517) );
  NOR4X1_LVT U637 ( .A1(n520), .A2(n519), .A3(n518), .A4(n517), .Y(n531) );
  AO22X1_LVT U638 ( .A1(n3462), .A2(\regs[18][17] ), .A3(n3476), .A4(
        \regs[14][17] ), .Y(n524) );
  AO22X1_LVT U639 ( .A1(n3465), .A2(\regs[10][17] ), .A3(n3489), .A4(
        \regs[22][17] ), .Y(n523) );
  AO22X1_LVT U640 ( .A1(n3454), .A2(\regs[2][17] ), .A3(n3484), .A4(
        \regs[27][17] ), .Y(n522) );
  AO22X1_LVT U641 ( .A1(n3485), .A2(\regs[8][17] ), .A3(n3490), .A4(
        \regs[11][17] ), .Y(n521) );
  NOR4X1_LVT U642 ( .A1(n524), .A2(n523), .A3(n522), .A4(n521), .Y(n530) );
  AO22X1_LVT U643 ( .A1(n3455), .A2(\regs[5][17] ), .A3(n3458), .A4(
        \regs[1][17] ), .Y(n528) );
  AO22X1_LVT U644 ( .A1(n3472), .A2(\regs[16][17] ), .A3(n3477), .A4(
        \regs[21][17] ), .Y(n527) );
  AO22X1_LVT U645 ( .A1(n3459), .A2(\regs[25][17] ), .A3(n3468), .A4(
        \regs[26][17] ), .Y(n526) );
  AO22X1_LVT U646 ( .A1(n3456), .A2(\regs[19][17] ), .A3(n3482), .A4(
        \regs[28][17] ), .Y(n525) );
  NOR4X1_LVT U647 ( .A1(n528), .A2(n527), .A3(n526), .A4(n525), .Y(n529) );
  NAND3X0_LVT U648 ( .A1(n531), .A2(n530), .A3(n529), .Y(n532) );
  OR3X1_LVT U649 ( .A1(n534), .A2(n533), .A3(n532), .Y(n535) );
  AO22X1_LVT U651 ( .A1(n8), .A2(n535), .A3(n79), .A4(wdata[17]), .Y(
        rdata2[17]) );
  AO22X1_LVT U652 ( .A1(n3490), .A2(\regs[11][18] ), .A3(n3477), .A4(
        \regs[21][18] ), .Y(n558) );
  AO22X1_LVT U653 ( .A1(n3473), .A2(\regs[30][18] ), .A3(n3476), .A4(
        \regs[14][18] ), .Y(n536) );
  INVX1_LVT U654 ( .A(n536), .Y(n540) );
  AO22X1_LVT U655 ( .A1(n3488), .A2(\regs[23][18] ), .A3(n3485), .A4(
        \regs[8][18] ), .Y(n537) );
  INVX1_LVT U656 ( .A(n537), .Y(n539) );
  NAND2X0_LVT U657 ( .A1(n3472), .A2(\regs[16][18] ), .Y(n538) );
  NAND3X0_LVT U658 ( .A1(n540), .A2(n539), .A3(n538), .Y(n557) );
  AO22X1_LVT U659 ( .A1(n3466), .A2(\regs[7][18] ), .A3(n3474), .A4(
        \regs[31][18] ), .Y(n544) );
  AO22X1_LVT U660 ( .A1(n3465), .A2(\regs[10][18] ), .A3(n3487), .A4(
        \regs[29][18] ), .Y(n543) );
  AO22X1_LVT U661 ( .A1(n3459), .A2(\regs[25][18] ), .A3(n3478), .A4(
        \regs[24][18] ), .Y(n542) );
  AO22X1_LVT U662 ( .A1(n3454), .A2(\regs[2][18] ), .A3(n3463), .A4(
        \regs[20][18] ), .Y(n541) );
  NOR4X1_LVT U663 ( .A1(n544), .A2(n543), .A3(n542), .A4(n541), .Y(n555) );
  AO22X1_LVT U664 ( .A1(n3460), .A2(\regs[4][18] ), .A3(n3489), .A4(
        \regs[22][18] ), .Y(n548) );
  AO22X1_LVT U665 ( .A1(n3484), .A2(\regs[27][18] ), .A3(n3464), .A4(
        \regs[13][18] ), .Y(n547) );
  AO22X1_LVT U666 ( .A1(n3462), .A2(\regs[18][18] ), .A3(n3482), .A4(
        \regs[28][18] ), .Y(n546) );
  AO22X1_LVT U667 ( .A1(n3479), .A2(\regs[6][18] ), .A3(n3467), .A4(
        \regs[17][18] ), .Y(n545) );
  NOR4X1_LVT U668 ( .A1(n548), .A2(n547), .A3(n546), .A4(n545), .Y(n554) );
  AO22X1_LVT U669 ( .A1(n3455), .A2(\regs[5][18] ), .A3(n3458), .A4(
        \regs[1][18] ), .Y(n552) );
  AO22X1_LVT U670 ( .A1(n3471), .A2(\regs[15][18] ), .A3(n3457), .A4(
        \regs[9][18] ), .Y(n551) );
  AO22X1_LVT U671 ( .A1(n3461), .A2(\regs[3][18] ), .A3(n3468), .A4(
        \regs[26][18] ), .Y(n550) );
  AO22X1_LVT U672 ( .A1(n3456), .A2(\regs[19][18] ), .A3(n3480), .A4(
        \regs[12][18] ), .Y(n549) );
  NOR4X1_LVT U673 ( .A1(n552), .A2(n551), .A3(n550), .A4(n549), .Y(n553) );
  NAND3X0_LVT U674 ( .A1(n555), .A2(n554), .A3(n553), .Y(n556) );
  OR3X1_LVT U675 ( .A1(n558), .A2(n557), .A3(n556), .Y(n559) );
  AO22X1_LVT U677 ( .A1(n8), .A2(n559), .A3(n79), .A4(n3491), .Y(rdata2[18])
         );
  AO22X1_LVT U678 ( .A1(n3473), .A2(\regs[30][19] ), .A3(n3484), .A4(
        \regs[27][19] ), .Y(n583) );
  AO22X1_LVT U679 ( .A1(n3476), .A2(\regs[14][19] ), .A3(n26), .A4(
        \regs[19][19] ), .Y(n560) );
  INVX1_LVT U680 ( .A(n560), .Y(n564) );
  AO22X1_LVT U681 ( .A1(n3460), .A2(\regs[4][19] ), .A3(n3488), .A4(
        \regs[23][19] ), .Y(n561) );
  INVX1_LVT U682 ( .A(n561), .Y(n563) );
  NAND2X0_LVT U683 ( .A1(n3462), .A2(\regs[18][19] ), .Y(n562) );
  NAND3X0_LVT U684 ( .A1(n564), .A2(n563), .A3(n562), .Y(n582) );
  AO22X1_LVT U685 ( .A1(n3466), .A2(\regs[7][19] ), .A3(n3489), .A4(
        \regs[22][19] ), .Y(n568) );
  AO22X1_LVT U686 ( .A1(n3463), .A2(\regs[20][19] ), .A3(n3477), .A4(
        \regs[21][19] ), .Y(n567) );
  AO22X1_LVT U687 ( .A1(n3457), .A2(\regs[9][19] ), .A3(n3474), .A4(
        \regs[31][19] ), .Y(n566) );
  AO22X1_LVT U688 ( .A1(n3465), .A2(\regs[10][19] ), .A3(n3458), .A4(
        \regs[1][19] ), .Y(n565) );
  NOR4X1_LVT U689 ( .A1(n568), .A2(n567), .A3(n566), .A4(n565), .Y(n580) );
  AO22X1_LVT U691 ( .A1(n3478), .A2(\regs[24][19] ), .A3(n3487), .A4(
        \regs[29][19] ), .Y(n573) );
  AO22X1_LVT U692 ( .A1(n3454), .A2(\regs[2][19] ), .A3(n3479), .A4(
        \regs[6][19] ), .Y(n572) );
  AO22X1_LVT U693 ( .A1(n3482), .A2(\regs[28][19] ), .A3(n3490), .A4(
        \regs[11][19] ), .Y(n571) );
  AO22X1_LVT U694 ( .A1(n3459), .A2(\regs[25][19] ), .A3(n3485), .A4(
        \regs[8][19] ), .Y(n570) );
  NOR4X1_LVT U695 ( .A1(n573), .A2(n572), .A3(n571), .A4(n570), .Y(n579) );
  AO22X1_LVT U696 ( .A1(n3455), .A2(\regs[5][19] ), .A3(n3464), .A4(
        \regs[13][19] ), .Y(n577) );
  AO22X1_LVT U697 ( .A1(n3461), .A2(\regs[3][19] ), .A3(n3468), .A4(
        \regs[26][19] ), .Y(n576) );
  AO22X1_LVT U698 ( .A1(n3472), .A2(\regs[16][19] ), .A3(n3480), .A4(
        \regs[12][19] ), .Y(n575) );
  AO22X1_LVT U699 ( .A1(n3471), .A2(\regs[15][19] ), .A3(n3467), .A4(
        \regs[17][19] ), .Y(n574) );
  NOR4X1_LVT U700 ( .A1(n577), .A2(n576), .A3(n575), .A4(n574), .Y(n578) );
  NAND3X0_LVT U701 ( .A1(n580), .A2(n579), .A3(n578), .Y(n581) );
  OR3X1_LVT U702 ( .A1(n583), .A2(n582), .A3(n581), .Y(n584) );
  AO22X1_LVT U704 ( .A1(n8), .A2(n584), .A3(n79), .A4(n3496), .Y(rdata2[19])
         );
  AO22X1_LVT U705 ( .A1(n3476), .A2(\regs[14][20] ), .A3(n3472), .A4(
        \regs[16][20] ), .Y(n607) );
  AO22X1_LVT U706 ( .A1(n3465), .A2(\regs[10][20] ), .A3(n3479), .A4(
        \regs[6][20] ), .Y(n585) );
  INVX1_LVT U707 ( .A(n585), .Y(n589) );
  AO22X1_LVT U708 ( .A1(n3458), .A2(\regs[1][20] ), .A3(n3457), .A4(
        \regs[9][20] ), .Y(n586) );
  INVX1_LVT U709 ( .A(n586), .Y(n588) );
  NAND2X0_LVT U710 ( .A1(n3464), .A2(\regs[13][20] ), .Y(n587) );
  NAND3X0_LVT U711 ( .A1(n589), .A2(n588), .A3(n587), .Y(n606) );
  AO22X1_LVT U712 ( .A1(n3456), .A2(\regs[19][20] ), .A3(n3478), .A4(
        \regs[24][20] ), .Y(n593) );
  AO22X1_LVT U713 ( .A1(n3460), .A2(\regs[4][20] ), .A3(n3482), .A4(
        \regs[28][20] ), .Y(n592) );
  AO22X1_LVT U714 ( .A1(n3471), .A2(\regs[15][20] ), .A3(n3468), .A4(
        \regs[26][20] ), .Y(n591) );
  AO22X1_LVT U715 ( .A1(n3473), .A2(\regs[30][20] ), .A3(n3490), .A4(
        \regs[11][20] ), .Y(n590) );
  NOR4X1_LVT U716 ( .A1(n593), .A2(n592), .A3(n591), .A4(n590), .Y(n604) );
  AO22X1_LVT U717 ( .A1(n3484), .A2(\regs[27][20] ), .A3(n3474), .A4(
        \regs[31][20] ), .Y(n597) );
  AO22X1_LVT U718 ( .A1(n3466), .A2(\regs[7][20] ), .A3(n3463), .A4(
        \regs[20][20] ), .Y(n596) );
  AO22X1_LVT U719 ( .A1(n3455), .A2(\regs[5][20] ), .A3(n3459), .A4(
        \regs[25][20] ), .Y(n595) );
  AO22X1_LVT U720 ( .A1(n3454), .A2(\regs[2][20] ), .A3(n3480), .A4(
        \regs[12][20] ), .Y(n594) );
  NOR4X1_LVT U721 ( .A1(n597), .A2(n596), .A3(n595), .A4(n594), .Y(n603) );
  AO22X1_LVT U722 ( .A1(n3489), .A2(\regs[22][20] ), .A3(n3467), .A4(
        \regs[17][20] ), .Y(n601) );
  AO22X1_LVT U723 ( .A1(n3461), .A2(\regs[3][20] ), .A3(n3488), .A4(
        \regs[23][20] ), .Y(n600) );
  AO22X1_LVT U724 ( .A1(n3462), .A2(\regs[18][20] ), .A3(n3485), .A4(
        \regs[8][20] ), .Y(n599) );
  AO22X1_LVT U725 ( .A1(n3477), .A2(\regs[21][20] ), .A3(n3487), .A4(
        \regs[29][20] ), .Y(n598) );
  NOR4X1_LVT U726 ( .A1(n601), .A2(n600), .A3(n599), .A4(n598), .Y(n602) );
  NAND3X0_LVT U727 ( .A1(n604), .A2(n603), .A3(n602), .Y(n605) );
  OR3X1_LVT U728 ( .A1(n607), .A2(n606), .A3(n605), .Y(n608) );
  AO22X1_LVT U730 ( .A1(n8), .A2(n608), .A3(n79), .A4(n3483), .Y(rdata2[20])
         );
  AO22X1_LVT U731 ( .A1(n3480), .A2(\regs[12][21] ), .A3(n3474), .A4(
        \regs[31][21] ), .Y(n632) );
  AO22X1_LVT U732 ( .A1(n3456), .A2(\regs[19][21] ), .A3(n3487), .A4(
        \regs[29][21] ), .Y(n609) );
  INVX1_LVT U733 ( .A(n609), .Y(n613) );
  AO22X1_LVT U734 ( .A1(n3460), .A2(\regs[4][21] ), .A3(n3463), .A4(
        \regs[20][21] ), .Y(n610) );
  INVX1_LVT U735 ( .A(n610), .Y(n612) );
  NAND2X0_LVT U736 ( .A1(n3490), .A2(\regs[11][21] ), .Y(n611) );
  NAND3X0_LVT U737 ( .A1(n613), .A2(n612), .A3(n611), .Y(n631) );
  AO22X1_LVT U738 ( .A1(n3476), .A2(\regs[14][21] ), .A3(n3457), .A4(
        \regs[9][21] ), .Y(n618) );
  AO22X1_LVT U739 ( .A1(n3466), .A2(\regs[7][21] ), .A3(n3479), .A4(
        \regs[6][21] ), .Y(n617) );
  AO22X1_LVT U740 ( .A1(n3473), .A2(\regs[30][21] ), .A3(n3484), .A4(
        \regs[27][21] ), .Y(n616) );
  AO22X1_LVT U741 ( .A1(n3464), .A2(\regs[13][21] ), .A3(n3472), .A4(
        \regs[16][21] ), .Y(n615) );
  NOR4X1_LVT U742 ( .A1(n618), .A2(n617), .A3(n616), .A4(n615), .Y(n629) );
  AO22X1_LVT U743 ( .A1(n3489), .A2(\regs[22][21] ), .A3(n3478), .A4(
        \regs[24][21] ), .Y(n622) );
  AO22X1_LVT U744 ( .A1(n3455), .A2(\regs[5][21] ), .A3(n3471), .A4(
        \regs[15][21] ), .Y(n621) );
  AO22X1_LVT U745 ( .A1(n3462), .A2(\regs[18][21] ), .A3(n3477), .A4(
        \regs[21][21] ), .Y(n620) );
  AO22X1_LVT U746 ( .A1(n3454), .A2(\regs[2][21] ), .A3(n3468), .A4(
        \regs[26][21] ), .Y(n619) );
  NOR4X1_LVT U747 ( .A1(n622), .A2(n621), .A3(n620), .A4(n619), .Y(n628) );
  AO22X1_LVT U748 ( .A1(n3459), .A2(\regs[25][21] ), .A3(n3488), .A4(
        \regs[23][21] ), .Y(n626) );
  AO22X1_LVT U749 ( .A1(n3482), .A2(\regs[28][21] ), .A3(n3461), .A4(
        \regs[3][21] ), .Y(n625) );
  AO22X1_LVT U750 ( .A1(n3485), .A2(\regs[8][21] ), .A3(n3467), .A4(
        \regs[17][21] ), .Y(n624) );
  AO22X1_LVT U751 ( .A1(n3465), .A2(\regs[10][21] ), .A3(n3458), .A4(
        \regs[1][21] ), .Y(n623) );
  NOR4X1_LVT U752 ( .A1(n626), .A2(n625), .A3(n624), .A4(n623), .Y(n627) );
  NAND3X0_LVT U753 ( .A1(n629), .A2(n628), .A3(n627), .Y(n630) );
  OR3X1_LVT U754 ( .A1(n632), .A2(n631), .A3(n630), .Y(n633) );
  AO22X1_LVT U756 ( .A1(n8), .A2(n633), .A3(n79), .A4(wdata[21]), .Y(
        rdata2[21]) );
  AO22X1_LVT U758 ( .A1(n3461), .A2(\regs[3][22] ), .A3(n3477), .A4(
        \regs[21][22] ), .Y(n662) );
  AO22X1_LVT U759 ( .A1(n3455), .A2(\regs[5][22] ), .A3(n3456), .A4(
        \regs[19][22] ), .Y(n636) );
  INVX1_LVT U760 ( .A(n636), .Y(n641) );
  AO22X1_LVT U761 ( .A1(n3462), .A2(\regs[18][22] ), .A3(n3474), .A4(
        \regs[31][22] ), .Y(n637) );
  INVX1_LVT U762 ( .A(n637), .Y(n640) );
  NAND2X0_LVT U763 ( .A1(n3487), .A2(\regs[29][22] ), .Y(n639) );
  NAND3X0_LVT U764 ( .A1(n641), .A2(n640), .A3(n639), .Y(n661) );
  AO22X1_LVT U766 ( .A1(n3484), .A2(\regs[27][22] ), .A3(n3479), .A4(
        \regs[6][22] ), .Y(n648) );
  AO22X1_LVT U767 ( .A1(n3465), .A2(\regs[10][22] ), .A3(n3472), .A4(
        \regs[16][22] ), .Y(n647) );
  AO22X1_LVT U768 ( .A1(n3466), .A2(\regs[7][22] ), .A3(n3490), .A4(
        \regs[11][22] ), .Y(n646) );
  AO22X1_LVT U769 ( .A1(n3478), .A2(\regs[24][22] ), .A3(n3467), .A4(
        \regs[17][22] ), .Y(n645) );
  NOR4X1_LVT U770 ( .A1(n648), .A2(n647), .A3(n646), .A4(n645), .Y(n659) );
  AO22X1_LVT U771 ( .A1(n3454), .A2(\regs[2][22] ), .A3(n3458), .A4(
        \regs[1][22] ), .Y(n652) );
  AO22X1_LVT U772 ( .A1(n3459), .A2(\regs[25][22] ), .A3(n3488), .A4(
        \regs[23][22] ), .Y(n651) );
  AO22X1_LVT U773 ( .A1(n3471), .A2(\regs[15][22] ), .A3(n3457), .A4(
        \regs[9][22] ), .Y(n650) );
  AO22X1_LVT U774 ( .A1(n3460), .A2(\regs[4][22] ), .A3(n3476), .A4(
        \regs[14][22] ), .Y(n649) );
  NOR4X1_LVT U775 ( .A1(n652), .A2(n651), .A3(n650), .A4(n649), .Y(n658) );
  AO22X1_LVT U776 ( .A1(n3464), .A2(\regs[13][22] ), .A3(n3485), .A4(
        \regs[8][22] ), .Y(n656) );
  AO22X1_LVT U777 ( .A1(n3489), .A2(\regs[22][22] ), .A3(n3480), .A4(
        \regs[12][22] ), .Y(n655) );
  AO22X1_LVT U778 ( .A1(n3473), .A2(\regs[30][22] ), .A3(n3468), .A4(
        \regs[26][22] ), .Y(n654) );
  AO22X1_LVT U779 ( .A1(n3482), .A2(\regs[28][22] ), .A3(n3463), .A4(
        \regs[20][22] ), .Y(n653) );
  NOR4X1_LVT U780 ( .A1(n656), .A2(n655), .A3(n654), .A4(n653), .Y(n657) );
  NAND3X0_LVT U781 ( .A1(n659), .A2(n658), .A3(n657), .Y(n660) );
  OR3X1_LVT U782 ( .A1(n662), .A2(n661), .A3(n660), .Y(n663) );
  AO22X1_LVT U784 ( .A1(n8), .A2(n663), .A3(n79), .A4(n3494), .Y(rdata2[22])
         );
  AO22X1_LVT U785 ( .A1(n3460), .A2(\regs[4][23] ), .A3(n3456), .A4(
        \regs[19][23] ), .Y(n688) );
  AO22X1_LVT U786 ( .A1(n3455), .A2(\regs[5][23] ), .A3(n3479), .A4(
        \regs[6][23] ), .Y(n664) );
  INVX1_LVT U787 ( .A(n664), .Y(n668) );
  AO22X1_LVT U788 ( .A1(n3465), .A2(\regs[10][23] ), .A3(n3457), .A4(
        \regs[9][23] ), .Y(n665) );
  INVX1_LVT U789 ( .A(n665), .Y(n667) );
  NAND2X0_LVT U790 ( .A1(n3458), .A2(\regs[1][23] ), .Y(n666) );
  NAND3X0_LVT U791 ( .A1(n668), .A2(n667), .A3(n666), .Y(n687) );
  AO22X1_LVT U792 ( .A1(n3454), .A2(\regs[2][23] ), .A3(n3489), .A4(
        \regs[22][23] ), .Y(n673) );
  AO22X1_LVT U793 ( .A1(n3474), .A2(\regs[31][23] ), .A3(n3487), .A4(
        \regs[29][23] ), .Y(n672) );
  AO22X1_LVT U794 ( .A1(n3471), .A2(\regs[15][23] ), .A3(n3462), .A4(
        \regs[18][23] ), .Y(n671) );
  AO22X1_LVT U795 ( .A1(n3464), .A2(\regs[13][23] ), .A3(n3485), .A4(
        \regs[8][23] ), .Y(n670) );
  NOR4X1_LVT U796 ( .A1(n673), .A2(n672), .A3(n671), .A4(n670), .Y(n685) );
  AO22X1_LVT U797 ( .A1(n3461), .A2(\regs[3][23] ), .A3(n3490), .A4(
        \regs[11][23] ), .Y(n678) );
  AO22X1_LVT U798 ( .A1(n3476), .A2(\regs[14][23] ), .A3(n40), .A4(
        \regs[20][23] ), .Y(n677) );
  AO22X1_LVT U799 ( .A1(n3472), .A2(\regs[16][23] ), .A3(n3480), .A4(
        \regs[12][23] ), .Y(n676) );
  AO22X1_LVT U801 ( .A1(n3468), .A2(\regs[26][23] ), .A3(n3477), .A4(
        \regs[21][23] ), .Y(n675) );
  NOR4X1_LVT U802 ( .A1(n678), .A2(n677), .A3(n676), .A4(n675), .Y(n684) );
  AO22X1_LVT U803 ( .A1(n3466), .A2(\regs[7][23] ), .A3(n3482), .A4(
        \regs[28][23] ), .Y(n682) );
  AO22X1_LVT U804 ( .A1(n3488), .A2(\regs[23][23] ), .A3(n3478), .A4(
        \regs[24][23] ), .Y(n681) );
  AO22X1_LVT U805 ( .A1(n3484), .A2(\regs[27][23] ), .A3(n3459), .A4(
        \regs[25][23] ), .Y(n680) );
  AO22X1_LVT U806 ( .A1(n3473), .A2(\regs[30][23] ), .A3(n3467), .A4(
        \regs[17][23] ), .Y(n679) );
  NOR4X1_LVT U807 ( .A1(n682), .A2(n681), .A3(n680), .A4(n679), .Y(n683) );
  NAND3X0_LVT U808 ( .A1(n685), .A2(n684), .A3(n683), .Y(n686) );
  OR3X1_LVT U809 ( .A1(n688), .A2(n687), .A3(n686), .Y(n689) );
  AO22X1_LVT U811 ( .A1(n8), .A2(n689), .A3(n79), .A4(n3497), .Y(rdata2[23])
         );
  AO22X1_LVT U812 ( .A1(n3459), .A2(\regs[25][24] ), .A3(n3457), .A4(
        \regs[9][24] ), .Y(n715) );
  AO22X1_LVT U813 ( .A1(n3465), .A2(\regs[10][24] ), .A3(n3488), .A4(
        \regs[23][24] ), .Y(n690) );
  INVX1_LVT U814 ( .A(n690), .Y(n695) );
  AO22X1_LVT U815 ( .A1(n3480), .A2(\regs[12][24] ), .A3(n3490), .A4(
        \regs[11][24] ), .Y(n692) );
  INVX1_LVT U816 ( .A(n692), .Y(n694) );
  NAND2X0_LVT U817 ( .A1(n3463), .A2(\regs[20][24] ), .Y(n693) );
  NAND3X0_LVT U818 ( .A1(n695), .A2(n694), .A3(n693), .Y(n714) );
  AO22X1_LVT U819 ( .A1(n3474), .A2(\regs[31][24] ), .A3(n3487), .A4(
        \regs[29][24] ), .Y(n701) );
  AO22X1_LVT U820 ( .A1(n3485), .A2(\regs[8][24] ), .A3(n3477), .A4(
        \regs[21][24] ), .Y(n700) );
  AO22X1_LVT U821 ( .A1(n3484), .A2(\regs[27][24] ), .A3(n3464), .A4(
        \regs[13][24] ), .Y(n699) );
  AO22X1_LVT U823 ( .A1(n3458), .A2(\regs[1][24] ), .A3(n3478), .A4(
        \regs[24][24] ), .Y(n698) );
  NOR4X1_LVT U824 ( .A1(n701), .A2(n700), .A3(n699), .A4(n698), .Y(n712) );
  AO22X1_LVT U825 ( .A1(n3454), .A2(\regs[2][24] ), .A3(n3479), .A4(
        \regs[6][24] ), .Y(n705) );
  AO22X1_LVT U826 ( .A1(n3472), .A2(\regs[16][24] ), .A3(n3468), .A4(
        \regs[26][24] ), .Y(n704) );
  AO22X1_LVT U827 ( .A1(n3466), .A2(\regs[7][24] ), .A3(n3456), .A4(
        \regs[19][24] ), .Y(n703) );
  AO22X1_LVT U828 ( .A1(n3462), .A2(\regs[18][24] ), .A3(n3489), .A4(
        \regs[22][24] ), .Y(n702) );
  NOR4X1_LVT U829 ( .A1(n705), .A2(n704), .A3(n703), .A4(n702), .Y(n711) );
  AO22X1_LVT U830 ( .A1(n3455), .A2(\regs[5][24] ), .A3(n3482), .A4(
        \regs[28][24] ), .Y(n709) );
  AO22X1_LVT U831 ( .A1(n3476), .A2(\regs[14][24] ), .A3(n3461), .A4(
        \regs[3][24] ), .Y(n708) );
  AO22X1_LVT U832 ( .A1(n3473), .A2(\regs[30][24] ), .A3(n3467), .A4(
        \regs[17][24] ), .Y(n707) );
  AO22X1_LVT U833 ( .A1(n3471), .A2(\regs[15][24] ), .A3(n3460), .A4(
        \regs[4][24] ), .Y(n706) );
  NOR4X1_LVT U834 ( .A1(n709), .A2(n708), .A3(n707), .A4(n706), .Y(n710) );
  NAND3X0_LVT U835 ( .A1(n712), .A2(n711), .A3(n710), .Y(n713) );
  OR3X1_LVT U836 ( .A1(n715), .A2(n714), .A3(n713), .Y(n716) );
  AO22X1_LVT U838 ( .A1(n8), .A2(n716), .A3(n79), .A4(n3493), .Y(rdata2[24])
         );
  AO22X1_LVT U839 ( .A1(n38), .A2(\regs[16][25] ), .A3(n39), .A4(
        \regs[23][25] ), .Y(n741) );
  AO22X1_LVT U840 ( .A1(n36), .A2(\regs[22][25] ), .A3(n61), .A4(
        \regs[24][25] ), .Y(n718) );
  INVX1_LVT U841 ( .A(n718), .Y(n722) );
  AO22X1_LVT U842 ( .A1(n21), .A2(\regs[30][25] ), .A3(n42), .A4(
        \regs[12][25] ), .Y(n719) );
  INVX1_LVT U843 ( .A(n719), .Y(n721) );
  NAND2X0_LVT U844 ( .A1(n25), .A2(\regs[14][25] ), .Y(n720) );
  NAND3X0_LVT U845 ( .A1(n722), .A2(n721), .A3(n720), .Y(n740) );
  AO22X1_LVT U846 ( .A1(n29), .A2(\regs[28][25] ), .A3(n3474), .A4(
        \regs[31][25] ), .Y(n726) );
  AO22X1_LVT U847 ( .A1(n37), .A2(\regs[3][25] ), .A3(n56), .A4(\regs[9][25] ), 
        .Y(n725) );
  AO22X1_LVT U848 ( .A1(n23), .A2(\regs[27][25] ), .A3(n63), .A4(
        \regs[17][25] ), .Y(n724) );
  AO22X1_LVT U849 ( .A1(n135), .A2(\regs[5][25] ), .A3(n54), .A4(
        \regs[21][25] ), .Y(n723) );
  NOR4X1_LVT U850 ( .A1(n726), .A2(n725), .A3(n724), .A4(n723), .Y(n738) );
  AO22X1_LVT U851 ( .A1(n3479), .A2(\regs[6][25] ), .A3(n40), .A4(
        \regs[20][25] ), .Y(n731) );
  AO22X1_LVT U852 ( .A1(n3466), .A2(\regs[7][25] ), .A3(n148), .A4(
        \regs[2][25] ), .Y(n730) );
  AO22X1_LVT U853 ( .A1(n30), .A2(\regs[25][25] ), .A3(n50), .A4(
        \regs[26][25] ), .Y(n729) );
  AO22X1_LVT U854 ( .A1(n3464), .A2(\regs[13][25] ), .A3(n65), .A4(
        \regs[29][25] ), .Y(n728) );
  NOR4X1_LVT U855 ( .A1(n731), .A2(n730), .A3(n729), .A4(n728), .Y(n737) );
  AO22X1_LVT U856 ( .A1(n110), .A2(\regs[18][25] ), .A3(n26), .A4(
        \regs[19][25] ), .Y(n735) );
  AO22X1_LVT U857 ( .A1(n43), .A2(\regs[8][25] ), .A3(n44), .A4(\regs[11][25] ), .Y(n734) );
  AO22X1_LVT U858 ( .A1(n120), .A2(\regs[4][25] ), .A3(n122), .A4(
        \regs[10][25] ), .Y(n733) );
  AO22X1_LVT U859 ( .A1(n3471), .A2(\regs[15][25] ), .A3(n52), .A4(
        \regs[1][25] ), .Y(n732) );
  NOR4X1_LVT U860 ( .A1(n735), .A2(n734), .A3(n733), .A4(n732), .Y(n736) );
  NAND3X0_LVT U861 ( .A1(n738), .A2(n737), .A3(n736), .Y(n739) );
  OR3X1_LVT U862 ( .A1(n741), .A2(n740), .A3(n739), .Y(n742) );
  AO22X1_LVT U864 ( .A1(n8), .A2(n742), .A3(n79), .A4(wdata[25]), .Y(
        rdata2[25]) );
  AO22X1_LVT U865 ( .A1(n135), .A2(\regs[5][26] ), .A3(n61), .A4(
        \regs[24][26] ), .Y(n765) );
  AO22X1_LVT U866 ( .A1(n3456), .A2(\regs[19][26] ), .A3(n3488), .A4(
        \regs[23][26] ), .Y(n743) );
  INVX1_LVT U867 ( .A(n743), .Y(n747) );
  AO22X1_LVT U868 ( .A1(n29), .A2(\regs[28][26] ), .A3(n36), .A4(
        \regs[22][26] ), .Y(n744) );
  INVX1_LVT U869 ( .A(n744), .Y(n746) );
  NAND2X0_LVT U870 ( .A1(n56), .A2(\regs[9][26] ), .Y(n745) );
  NAND3X0_LVT U871 ( .A1(n747), .A2(n746), .A3(n745), .Y(n764) );
  AO22X1_LVT U872 ( .A1(n54), .A2(\regs[21][26] ), .A3(n58), .A4(
        \regs[31][26] ), .Y(n751) );
  AO22X1_LVT U873 ( .A1(n21), .A2(\regs[30][26] ), .A3(n42), .A4(
        \regs[12][26] ), .Y(n750) );
  AO22X1_LVT U874 ( .A1(n148), .A2(\regs[2][26] ), .A3(n3459), .A4(
        \regs[25][26] ), .Y(n749) );
  AO22X1_LVT U875 ( .A1(n9), .A2(\regs[15][26] ), .A3(n44), .A4(\regs[11][26] ), .Y(n748) );
  NOR4X1_LVT U876 ( .A1(n751), .A2(n750), .A3(n749), .A4(n748), .Y(n762) );
  AO22X1_LVT U877 ( .A1(n25), .A2(\regs[14][26] ), .A3(n65), .A4(
        \regs[29][26] ), .Y(n755) );
  AO22X1_LVT U878 ( .A1(n23), .A2(\regs[27][26] ), .A3(n37), .A4(\regs[3][26] ), .Y(n754) );
  AO22X1_LVT U879 ( .A1(n11), .A2(\regs[7][26] ), .A3(n63), .A4(\regs[17][26] ), .Y(n753) );
  AO22X1_LVT U880 ( .A1(n24), .A2(\regs[13][26] ), .A3(n43), .A4(\regs[8][26] ), .Y(n752) );
  NOR4X1_LVT U881 ( .A1(n755), .A2(n754), .A3(n753), .A4(n752), .Y(n761) );
  AO22X1_LVT U882 ( .A1(n122), .A2(\regs[10][26] ), .A3(n38), .A4(
        \regs[16][26] ), .Y(n759) );
  AO22X1_LVT U883 ( .A1(n120), .A2(\regs[4][26] ), .A3(n28), .A4(\regs[6][26] ), .Y(n758) );
  AO22X1_LVT U884 ( .A1(n110), .A2(\regs[18][26] ), .A3(n50), .A4(
        \regs[26][26] ), .Y(n757) );
  AO22X1_LVT U885 ( .A1(n40), .A2(\regs[20][26] ), .A3(n52), .A4(\regs[1][26] ), .Y(n756) );
  NOR4X1_LVT U886 ( .A1(n759), .A2(n758), .A3(n757), .A4(n756), .Y(n760) );
  NAND3X0_LVT U887 ( .A1(n762), .A2(n761), .A3(n760), .Y(n763) );
  OR3X1_LVT U888 ( .A1(n765), .A2(n764), .A3(n763), .Y(n766) );
  AO22X1_LVT U890 ( .A1(n8), .A2(n766), .A3(n79), .A4(n3503), .Y(rdata2[26])
         );
  AO22X1_LVT U891 ( .A1(n40), .A2(\regs[20][27] ), .A3(n3467), .A4(
        \regs[17][27] ), .Y(n790) );
  AO22X1_LVT U892 ( .A1(n39), .A2(\regs[23][27] ), .A3(n3457), .A4(
        \regs[9][27] ), .Y(n767) );
  INVX1_LVT U893 ( .A(n767), .Y(n772) );
  AO22X1_LVT U894 ( .A1(n37), .A2(\regs[3][27] ), .A3(n38), .A4(\regs[16][27] ), .Y(n768) );
  INVX1_LVT U895 ( .A(n768), .Y(n771) );
  NAND2X0_LVT U896 ( .A1(n26), .A2(\regs[19][27] ), .Y(n770) );
  NAND3X0_LVT U897 ( .A1(n772), .A2(n771), .A3(n770), .Y(n789) );
  AO22X1_LVT U898 ( .A1(n9), .A2(\regs[15][27] ), .A3(n24), .A4(\regs[13][27] ), .Y(n776) );
  AO22X1_LVT U899 ( .A1(n23), .A2(\regs[27][27] ), .A3(n28), .A4(\regs[6][27] ), .Y(n775) );
  AO22X1_LVT U900 ( .A1(n3482), .A2(\regs[28][27] ), .A3(n3458), .A4(
        \regs[1][27] ), .Y(n774) );
  AO22X1_LVT U901 ( .A1(n21), .A2(\regs[30][27] ), .A3(n42), .A4(
        \regs[12][27] ), .Y(n773) );
  NOR4X1_LVT U902 ( .A1(n776), .A2(n775), .A3(n774), .A4(n773), .Y(n787) );
  AO22X1_LVT U903 ( .A1(n135), .A2(\regs[5][27] ), .A3(n36), .A4(
        \regs[22][27] ), .Y(n780) );
  AO22X1_LVT U904 ( .A1(n148), .A2(\regs[2][27] ), .A3(n3490), .A4(
        \regs[11][27] ), .Y(n779) );
  AO22X1_LVT U905 ( .A1(n58), .A2(\regs[31][27] ), .A3(n61), .A4(
        \regs[24][27] ), .Y(n778) );
  AO22X1_LVT U906 ( .A1(n3460), .A2(\regs[4][27] ), .A3(n50), .A4(
        \regs[26][27] ), .Y(n777) );
  NOR4X1_LVT U907 ( .A1(n780), .A2(n779), .A3(n778), .A4(n777), .Y(n786) );
  AO22X1_LVT U908 ( .A1(n30), .A2(\regs[25][27] ), .A3(n43), .A4(\regs[8][27] ), .Y(n784) );
  AO22X1_LVT U909 ( .A1(n3477), .A2(\regs[21][27] ), .A3(n65), .A4(
        \regs[29][27] ), .Y(n783) );
  AO22X1_LVT U910 ( .A1(n110), .A2(\regs[18][27] ), .A3(n3476), .A4(
        \regs[14][27] ), .Y(n782) );
  AO22X1_LVT U911 ( .A1(n122), .A2(\regs[10][27] ), .A3(n11), .A4(
        \regs[7][27] ), .Y(n781) );
  NOR4X1_LVT U912 ( .A1(n784), .A2(n783), .A3(n782), .A4(n781), .Y(n785) );
  NAND3X0_LVT U913 ( .A1(n787), .A2(n786), .A3(n785), .Y(n788) );
  OR3X1_LVT U914 ( .A1(n790), .A2(n789), .A3(n788), .Y(n791) );
  AO22X1_LVT U916 ( .A1(n8), .A2(n791), .A3(n79), .A4(wdata[27]), .Y(
        rdata2[27]) );
  AO22X1_LVT U917 ( .A1(n58), .A2(\regs[31][28] ), .A3(n61), .A4(
        \regs[24][28] ), .Y(n817) );
  AO22X1_LVT U918 ( .A1(n40), .A2(\regs[20][28] ), .A3(n65), .A4(
        \regs[29][28] ), .Y(n794) );
  INVX1_LVT U919 ( .A(n794), .Y(n798) );
  AO22X1_LVT U920 ( .A1(n11), .A2(\regs[7][28] ), .A3(n28), .A4(\regs[6][28] ), 
        .Y(n795) );
  INVX1_LVT U921 ( .A(n795), .Y(n797) );
  NAND2X0_LVT U922 ( .A1(n120), .A2(\regs[4][28] ), .Y(n796) );
  NAND3X0_LVT U923 ( .A1(n798), .A2(n797), .A3(n796), .Y(n816) );
  AO22X1_LVT U924 ( .A1(n29), .A2(\regs[28][28] ), .A3(n52), .A4(\regs[1][28] ), .Y(n802) );
  AO22X1_LVT U925 ( .A1(n23), .A2(\regs[27][28] ), .A3(n30), .A4(
        \regs[25][28] ), .Y(n801) );
  AO22X1_LVT U926 ( .A1(n148), .A2(\regs[2][28] ), .A3(n38), .A4(
        \regs[16][28] ), .Y(n800) );
  AO22X1_LVT U927 ( .A1(n26), .A2(\regs[19][28] ), .A3(n63), .A4(
        \regs[17][28] ), .Y(n799) );
  NOR4X1_LVT U928 ( .A1(n802), .A2(n801), .A3(n800), .A4(n799), .Y(n814) );
  AO22X1_LVT U929 ( .A1(n122), .A2(\regs[10][28] ), .A3(n56), .A4(
        \regs[9][28] ), .Y(n807) );
  AO22X1_LVT U930 ( .A1(n36), .A2(\regs[22][28] ), .A3(n44), .A4(
        \regs[11][28] ), .Y(n806) );
  AO22X1_LVT U931 ( .A1(n110), .A2(\regs[18][28] ), .A3(n21), .A4(
        \regs[30][28] ), .Y(n805) );
  AO22X1_LVT U932 ( .A1(n37), .A2(\regs[3][28] ), .A3(n39), .A4(\regs[23][28] ), .Y(n804) );
  NOR4X1_LVT U933 ( .A1(n807), .A2(n806), .A3(n805), .A4(n804), .Y(n813) );
  AO22X1_LVT U934 ( .A1(n50), .A2(\regs[26][28] ), .A3(n54), .A4(
        \regs[21][28] ), .Y(n811) );
  AO22X1_LVT U935 ( .A1(n24), .A2(\regs[13][28] ), .A3(n25), .A4(
        \regs[14][28] ), .Y(n810) );
  AO22X1_LVT U936 ( .A1(n135), .A2(\regs[5][28] ), .A3(n43), .A4(\regs[8][28] ), .Y(n809) );
  AO22X1_LVT U937 ( .A1(n9), .A2(\regs[15][28] ), .A3(n42), .A4(\regs[12][28] ), .Y(n808) );
  NOR4X1_LVT U938 ( .A1(n811), .A2(n810), .A3(n809), .A4(n808), .Y(n812) );
  NAND3X0_LVT U939 ( .A1(n814), .A2(n813), .A3(n812), .Y(n815) );
  OR3X1_LVT U940 ( .A1(n817), .A2(n816), .A3(n815), .Y(n818) );
  AO22X1_LVT U942 ( .A1(n8), .A2(n818), .A3(n79), .A4(n3500), .Y(rdata2[28])
         );
  AO22X1_LVT U943 ( .A1(n3456), .A2(\regs[19][29] ), .A3(n3489), .A4(
        \regs[22][29] ), .Y(n846) );
  AO22X1_LVT U944 ( .A1(n3485), .A2(\regs[8][29] ), .A3(n52), .A4(
        \regs[1][29] ), .Y(n820) );
  INVX1_LVT U945 ( .A(n820), .Y(n825) );
  AO22X1_LVT U946 ( .A1(n21), .A2(\regs[30][29] ), .A3(n42), .A4(
        \regs[12][29] ), .Y(n821) );
  INVX1_LVT U947 ( .A(n821), .Y(n824) );
  NAND2X0_LVT U948 ( .A1(n44), .A2(\regs[11][29] ), .Y(n823) );
  NAND3X0_LVT U949 ( .A1(n825), .A2(n824), .A3(n823), .Y(n845) );
  AO22X1_LVT U950 ( .A1(n135), .A2(\regs[5][29] ), .A3(n24), .A4(
        \regs[13][29] ), .Y(n830) );
  AO22X1_LVT U951 ( .A1(n3468), .A2(\regs[26][29] ), .A3(n65), .A4(
        \regs[29][29] ), .Y(n829) );
  AO22X1_LVT U952 ( .A1(n3460), .A2(\regs[4][29] ), .A3(n40), .A4(
        \regs[20][29] ), .Y(n828) );
  AO22X1_LVT U953 ( .A1(n39), .A2(\regs[23][29] ), .A3(n63), .A4(
        \regs[17][29] ), .Y(n827) );
  NOR4X1_LVT U954 ( .A1(n830), .A2(n829), .A3(n828), .A4(n827), .Y(n843) );
  AO22X1_LVT U955 ( .A1(n25), .A2(\regs[14][29] ), .A3(n38), .A4(
        \regs[16][29] ), .Y(n836) );
  AO22X1_LVT U956 ( .A1(n30), .A2(\regs[25][29] ), .A3(n37), .A4(\regs[3][29] ), .Y(n835) );
  AO22X1_LVT U957 ( .A1(n23), .A2(\regs[27][29] ), .A3(n54), .A4(
        \regs[21][29] ), .Y(n834) );
  AO22X1_LVT U958 ( .A1(n11), .A2(\regs[7][29] ), .A3(n28), .A4(\regs[6][29] ), 
        .Y(n833) );
  NOR4X1_LVT U959 ( .A1(n836), .A2(n835), .A3(n834), .A4(n833), .Y(n842) );
  AO22X1_LVT U960 ( .A1(n122), .A2(\regs[10][29] ), .A3(n56), .A4(
        \regs[9][29] ), .Y(n840) );
  AO22X1_LVT U961 ( .A1(n148), .A2(\regs[2][29] ), .A3(n3478), .A4(
        \regs[24][29] ), .Y(n839) );
  AO22X1_LVT U962 ( .A1(n9), .A2(\regs[15][29] ), .A3(n29), .A4(\regs[28][29] ), .Y(n838) );
  AO22X1_LVT U963 ( .A1(n110), .A2(\regs[18][29] ), .A3(n58), .A4(
        \regs[31][29] ), .Y(n837) );
  NOR4X1_LVT U964 ( .A1(n840), .A2(n839), .A3(n838), .A4(n837), .Y(n841) );
  NAND3X0_LVT U965 ( .A1(n843), .A2(n842), .A3(n841), .Y(n844) );
  OR3X1_LVT U966 ( .A1(n846), .A2(n845), .A3(n844), .Y(n848) );
  AO22X1_LVT U968 ( .A1(n8), .A2(n848), .A3(n79), .A4(n3501), .Y(rdata2[29])
         );
  AO22X1_LVT U970 ( .A1(n3454), .A2(\regs[2][30] ), .A3(n3463), .A4(
        \regs[20][30] ), .Y(n892) );
  AO22X1_LVT U971 ( .A1(n23), .A2(\regs[27][30] ), .A3(n58), .A4(
        \regs[31][30] ), .Y(n852) );
  INVX1_LVT U972 ( .A(n852), .Y(n859) );
  AO22X1_LVT U973 ( .A1(n24), .A2(\regs[13][30] ), .A3(n30), .A4(
        \regs[25][30] ), .Y(n855) );
  INVX1_LVT U974 ( .A(n855), .Y(n858) );
  NAND2X0_LVT U975 ( .A1(n54), .A2(\regs[21][30] ), .Y(n857) );
  NAND3X0_LVT U976 ( .A1(n859), .A2(n858), .A3(n857), .Y(n891) );
  AO22X1_LVT U977 ( .A1(n122), .A2(\regs[10][30] ), .A3(n42), .A4(
        \regs[12][30] ), .Y(n868) );
  AO22X1_LVT U978 ( .A1(n120), .A2(\regs[4][30] ), .A3(n28), .A4(\regs[6][30] ), .Y(n867) );
  AO22X1_LVT U979 ( .A1(n29), .A2(\regs[28][30] ), .A3(n65), .A4(
        \regs[29][30] ), .Y(n866) );
  AO22X1_LVT U980 ( .A1(n39), .A2(\regs[23][30] ), .A3(n44), .A4(
        \regs[11][30] ), .Y(n865) );
  NOR4X1_LVT U981 ( .A1(n868), .A2(n867), .A3(n866), .A4(n865), .Y(n889) );
  AO22X1_LVT U982 ( .A1(n11), .A2(\regs[7][30] ), .A3(n56), .A4(\regs[9][30] ), 
        .Y(n877) );
  AO22X1_LVT U983 ( .A1(n37), .A2(\regs[3][30] ), .A3(n38), .A4(\regs[16][30] ), .Y(n876) );
  AO22X1_LVT U984 ( .A1(n26), .A2(\regs[19][30] ), .A3(n36), .A4(
        \regs[22][30] ), .Y(n875) );
  AO22X1_LVT U985 ( .A1(n43), .A2(\regs[8][30] ), .A3(n50), .A4(\regs[26][30] ), .Y(n874) );
  NOR4X1_LVT U986 ( .A1(n877), .A2(n876), .A3(n875), .A4(n874), .Y(n888) );
  AO22X1_LVT U987 ( .A1(n21), .A2(\regs[30][30] ), .A3(n25), .A4(
        \regs[14][30] ), .Y(n886) );
  AO22X1_LVT U988 ( .A1(n9), .A2(\regs[15][30] ), .A3(n63), .A4(\regs[17][30] ), .Y(n885) );
  AO22X1_LVT U989 ( .A1(n135), .A2(\regs[5][30] ), .A3(n61), .A4(
        \regs[24][30] ), .Y(n884) );
  AO22X1_LVT U990 ( .A1(n3462), .A2(\regs[18][30] ), .A3(n3458), .A4(
        \regs[1][30] ), .Y(n883) );
  NOR4X1_LVT U991 ( .A1(n886), .A2(n885), .A3(n884), .A4(n883), .Y(n887) );
  NAND3X0_LVT U992 ( .A1(n889), .A2(n888), .A3(n887), .Y(n890) );
  OR3X1_LVT U993 ( .A1(n892), .A2(n891), .A3(n890), .Y(n894) );
  AO22X1_LVT U996 ( .A1(n8), .A2(n894), .A3(n79), .A4(wdata[30]), .Y(
        rdata2[30]) );
  AO22X1_LVT U997 ( .A1(n120), .A2(\regs[4][31] ), .A3(n63), .A4(
        \regs[17][31] ), .Y(n948) );
  AO22X1_LVT U998 ( .A1(n135), .A2(\regs[5][31] ), .A3(n9), .A4(\regs[15][31] ), .Y(n899) );
  INVX1_LVT U999 ( .A(n899), .Y(n906) );
  AO22X1_LVT U1000 ( .A1(n29), .A2(\regs[28][31] ), .A3(n3480), .A4(
        \regs[12][31] ), .Y(n902) );
  INVX1_LVT U1001 ( .A(n902), .Y(n905) );
  NAND2X0_LVT U1002 ( .A1(n50), .A2(\regs[26][31] ), .Y(n904) );
  NAND3X0_LVT U1003 ( .A1(n906), .A2(n905), .A3(n904), .Y(n947) );
  AO22X1_LVT U1004 ( .A1(n36), .A2(\regs[22][31] ), .A3(n3472), .A4(
        \regs[16][31] ), .Y(n918) );
  AO22X1_LVT U1005 ( .A1(n24), .A2(\regs[13][31] ), .A3(n54), .A4(
        \regs[21][31] ), .Y(n917) );
  AO22X1_LVT U1006 ( .A1(n11), .A2(\regs[7][31] ), .A3(n40), .A4(
        \regs[20][31] ), .Y(n916) );
  AO22X1_LVT U1007 ( .A1(n23), .A2(\regs[27][31] ), .A3(n58), .A4(
        \regs[31][31] ), .Y(n915) );
  NOR4X1_LVT U1008 ( .A1(n918), .A2(n917), .A3(n916), .A4(n915), .Y(n945) );
  AO22X1_LVT U1009 ( .A1(n122), .A2(\regs[10][31] ), .A3(n43), .A4(
        \regs[8][31] ), .Y(n930) );
  AO22X1_LVT U1010 ( .A1(n148), .A2(\regs[2][31] ), .A3(n44), .A4(
        \regs[11][31] ), .Y(n929) );
  AO22X1_LVT U1011 ( .A1(n21), .A2(\regs[30][31] ), .A3(n25), .A4(
        \regs[14][31] ), .Y(n928) );
  AO22X1_LVT U1012 ( .A1(n37), .A2(\regs[3][31] ), .A3(n39), .A4(
        \regs[23][31] ), .Y(n927) );
  NOR4X1_LVT U1013 ( .A1(n930), .A2(n929), .A3(n928), .A4(n927), .Y(n944) );
  AO22X1_LVT U1014 ( .A1(n26), .A2(\regs[19][31] ), .A3(n3479), .A4(
        \regs[6][31] ), .Y(n942) );
  AO22X1_LVT U1015 ( .A1(n52), .A2(\regs[1][31] ), .A3(n61), .A4(
        \regs[24][31] ), .Y(n941) );
  AO22X1_LVT U1016 ( .A1(n110), .A2(\regs[18][31] ), .A3(n65), .A4(
        \regs[29][31] ), .Y(n940) );
  AO22X1_LVT U1017 ( .A1(n30), .A2(\regs[25][31] ), .A3(n56), .A4(
        \regs[9][31] ), .Y(n939) );
  NOR4X1_LVT U1018 ( .A1(n942), .A2(n941), .A3(n940), .A4(n939), .Y(n943) );
  NAND3X0_LVT U1019 ( .A1(n945), .A2(n944), .A3(n943), .Y(n946) );
  OR3X1_LVT U1020 ( .A1(n948), .A2(n947), .A3(n946), .Y(n950) );
  AO22X1_LVT U1022 ( .A1(n8), .A2(n950), .A3(n79), .A4(n3486), .Y(rdata2[31])
         );
  OA22X1_LVT U1026 ( .A1(waddr[4]), .A2(n3452), .A3(waddr[3]), .A4(n3451), .Y(
        n952) );
  OA221X1_LVT U1027 ( .A1(n3077), .A2(raddr1[3]), .A3(n3002), .A4(raddr1[4]), 
        .A5(n952), .Y(n956) );
  INVX1_LVT U1028 ( .A(raddr1[0]), .Y(n971) );
  INVX1_LVT U1029 ( .A(raddr1[1]), .Y(n966) );
  OA22X1_LVT U1030 ( .A1(waddr[0]), .A2(n971), .A3(waddr[1]), .A4(n966), .Y(
        n953) );
  OA221X1_LVT U1031 ( .A1(n3192), .A2(raddr1[1]), .A3(n3191), .A4(raddr1[0]), 
        .A5(n953), .Y(n955) );
  AO22X1_LVT U1033 ( .A1(waddr[2]), .A2(raddr1[2]), .A3(n3298), .A4(n3450), 
        .Y(n954) );
  NAND4X0_LVT U1034 ( .A1(we), .A2(n956), .A3(n955), .A4(n954), .Y(n961) );
  INVX1_LVT U1035 ( .A(n961), .Y(n959) );
  AND2X1_LVT U1036 ( .A1(n3297), .A2(re1), .Y(n958) );
  NAND2X0_LVT U1037 ( .A1(n971), .A2(n966), .Y(n980) );
  NAND3X0_LVT U1038 ( .A1(n3450), .A2(n3452), .A3(n3451), .Y(n964) );
  OR2X1_LVT U1039 ( .A1(n980), .A2(n964), .Y(n957) );
  AND2X1_LVT U1040 ( .A1(n958), .A2(n957), .Y(n962) );
  INVX1_LVT U1047 ( .A(n964), .Y(n1013) );
  AND2X1_LVT U1048 ( .A1(raddr1[0]), .A2(raddr1[1]), .Y(n1026) );
  AND2X1_LVT U1052 ( .A1(raddr1[0]), .A2(n966), .Y(n1024) );
  AND3X1_LVT U1053 ( .A1(raddr1[3]), .A2(n3450), .A3(n3452), .Y(n1021) );
  AO22X1_LVT U1057 ( .A1(\regs[3][0] ), .A2(n965), .A3(\regs[9][0] ), .A4(n967), .Y(n1037) );
  AND3X1_LVT U1058 ( .A1(raddr1[4]), .A2(raddr1[2]), .A3(n3451), .Y(n1000) );
  AO22X1_LVT U1065 ( .A1(\regs[23][0] ), .A2(n968), .A3(\regs[21][0] ), .A4(
        n969), .Y(n970) );
  INVX1_LVT U1066 ( .A(n970), .Y(n978) );
  AND2X1_LVT U1067 ( .A1(raddr1[1]), .A2(n971), .Y(n1019) );
  AO22X1_LVT U1074 ( .A1(\regs[10][0] ), .A2(n972), .A3(\regs[29][0] ), .A4(
        n973), .Y(n974) );
  INVX1_LVT U1075 ( .A(n974), .Y(n977) );
  NAND2X0_LVT U1079 ( .A1(\regs[30][0] ), .A2(n975), .Y(n976) );
  NAND3X0_LVT U1080 ( .A1(n978), .A2(n977), .A3(n976), .Y(n1036) );
  AND3X1_LVT U1081 ( .A1(raddr1[4]), .A2(raddr1[3]), .A3(n3450), .Y(n1004) );
  INVX1_LVT U1085 ( .A(n980), .Y(n1011) );
  AO22X1_LVT U1089 ( .A1(\regs[25][0] ), .A2(n979), .A3(\regs[8][0] ), .A4(
        n981), .Y(n994) );
  AND3X1_LVT U1093 ( .A1(raddr1[2]), .A2(raddr1[3]), .A3(n3452), .Y(n1023) );
  AO22X1_LVT U1097 ( .A1(\regs[27][0] ), .A2(n982), .A3(\regs[12][0] ), .A4(
        n983), .Y(n993) );
  AND3X1_LVT U1098 ( .A1(raddr1[2]), .A2(n3452), .A3(n3451), .Y(n1018) );
  AO22X1_LVT U1105 ( .A1(\regs[7][0] ), .A2(n985), .A3(\regs[28][0] ), .A4(
        n986), .Y(n992) );
  AND3X1_LVT U1109 ( .A1(raddr1[4]), .A2(n3450), .A3(n3451), .Y(n1016) );
  AO22X1_LVT U1113 ( .A1(\regs[5][0] ), .A2(n987), .A3(\regs[17][0] ), .A4(
        n990), .Y(n991) );
  NOR4X1_LVT U1114 ( .A1(n994), .A2(n993), .A3(n992), .A4(n991), .Y(n1034) );
  AO22X1_LVT U1121 ( .A1(\regs[18][0] ), .A2(n995), .A3(\regs[22][0] ), .A4(
        n996), .Y(n1010) );
  AO22X1_LVT U1128 ( .A1(\regs[14][0] ), .A2(n997), .A3(\regs[1][0] ), .A4(
        n998), .Y(n1009) );
  AO22X1_LVT U1135 ( .A1(\regs[20][0] ), .A2(n1001), .A3(\regs[26][0] ), .A4(
        n1002), .Y(n1008) );
  AO22X1_LVT U1142 ( .A1(\regs[16][0] ), .A2(n1003), .A3(\regs[24][0] ), .A4(
        n1005), .Y(n1007) );
  NOR4X1_LVT U1143 ( .A1(n1010), .A2(n1009), .A3(n1008), .A4(n1007), .Y(n1033)
         );
  AO22X1_LVT U1150 ( .A1(\regs[4][0] ), .A2(n1012), .A3(\regs[2][0] ), .A4(
        n1014), .Y(n1031) );
  AO22X1_LVT U1157 ( .A1(\regs[15][0] ), .A2(n1015), .A3(\regs[19][0] ), .A4(
        n1017), .Y(n1030) );
  AO22X1_LVT U1164 ( .A1(\regs[6][0] ), .A2(n1020), .A3(\regs[11][0] ), .A4(
        n1022), .Y(n1029) );
  AO22X1_LVT U1171 ( .A1(\regs[13][0] ), .A2(n1025), .A3(\regs[31][0] ), .A4(
        n1027), .Y(n1028) );
  NOR4X1_LVT U1172 ( .A1(n1031), .A2(n1030), .A3(n1029), .A4(n1028), .Y(n1032)
         );
  NAND3X0_LVT U1173 ( .A1(n1034), .A2(n1033), .A3(n1032), .Y(n1035) );
  OR3X1_LVT U1174 ( .A1(n1037), .A2(n1036), .A3(n1035), .Y(n1038) );
  AO22X1_LVT U1175 ( .A1(wdata[0]), .A2(n960), .A3(n963), .A4(n1038), .Y(
        rdata1[0]) );
  AO22X1_LVT U1179 ( .A1(\regs[15][1] ), .A2(n1015), .A3(\regs[13][1] ), .A4(
        n1025), .Y(n1067) );
  AO22X1_LVT U1180 ( .A1(\regs[20][1] ), .A2(n1001), .A3(\regs[8][1] ), .A4(
        n981), .Y(n1040) );
  INVX1_LVT U1181 ( .A(n1040), .Y(n1045) );
  AO22X1_LVT U1183 ( .A1(\regs[1][1] ), .A2(n998), .A3(\regs[22][1] ), .A4(
        n996), .Y(n1042) );
  INVX1_LVT U1184 ( .A(n1042), .Y(n1044) );
  NAND2X0_LVT U1186 ( .A1(\regs[14][1] ), .A2(n997), .Y(n1043) );
  NAND3X0_LVT U1187 ( .A1(n1045), .A2(n1044), .A3(n1043), .Y(n1066) );
  AO22X1_LVT U1189 ( .A1(\regs[2][1] ), .A2(n1014), .A3(\regs[16][1] ), .A4(
        n1003), .Y(n1051) );
  AO22X1_LVT U1191 ( .A1(\regs[19][1] ), .A2(n1017), .A3(\regs[28][1] ), .A4(
        n986), .Y(n1050) );
  AO22X1_LVT U1194 ( .A1(\regs[12][1] ), .A2(n983), .A3(\regs[7][1] ), .A4(
        n985), .Y(n1049) );
  AO22X1_LVT U1197 ( .A1(\regs[5][1] ), .A2(n987), .A3(\regs[10][1] ), .A4(
        n972), .Y(n1048) );
  NOR4X1_LVT U1198 ( .A1(n1051), .A2(n1050), .A3(n1049), .A4(n1048), .Y(n1064)
         );
  AO22X1_LVT U1201 ( .A1(\regs[24][1] ), .A2(n1005), .A3(\regs[3][1] ), .A4(
        n965), .Y(n1057) );
  AO22X1_LVT U1204 ( .A1(\regs[9][1] ), .A2(n967), .A3(\regs[29][1] ), .A4(
        n973), .Y(n1056) );
  AO22X1_LVT U1207 ( .A1(\regs[21][1] ), .A2(n969), .A3(\regs[31][1] ), .A4(
        n1027), .Y(n1055) );
  AO22X1_LVT U1209 ( .A1(\regs[11][1] ), .A2(n1022), .A3(\regs[23][1] ), .A4(
        n968), .Y(n1054) );
  NOR4X1_LVT U1210 ( .A1(n1057), .A2(n1056), .A3(n1055), .A4(n1054), .Y(n1063)
         );
  AO22X1_LVT U1212 ( .A1(\regs[27][1] ), .A2(n982), .A3(\regs[4][1] ), .A4(
        n1012), .Y(n1061) );
  AO22X1_LVT U1215 ( .A1(\regs[30][1] ), .A2(n975), .A3(\regs[6][1] ), .A4(
        n1020), .Y(n1060) );
  AO22X1_LVT U1218 ( .A1(\regs[26][1] ), .A2(n1002), .A3(\regs[25][1] ), .A4(
        n979), .Y(n1059) );
  AO22X1_LVT U1220 ( .A1(\regs[18][1] ), .A2(n995), .A3(\regs[17][1] ), .A4(
        n990), .Y(n1058) );
  NOR4X1_LVT U1221 ( .A1(n1061), .A2(n1060), .A3(n1059), .A4(n1058), .Y(n1062)
         );
  NAND3X0_LVT U1222 ( .A1(n1064), .A2(n1063), .A3(n1062), .Y(n1065) );
  OR3X1_LVT U1223 ( .A1(n1067), .A2(n1066), .A3(n1065), .Y(n1068) );
  AO22X1_LVT U1224 ( .A1(wdata[1]), .A2(n960), .A3(n963), .A4(n1068), .Y(
        rdata1[1]) );
  AO22X1_LVT U1227 ( .A1(\regs[7][2] ), .A2(n985), .A3(\regs[5][2] ), .A4(n987), .Y(n1106) );
  AO22X1_LVT U1230 ( .A1(\regs[22][2] ), .A2(n996), .A3(\regs[30][2] ), .A4(
        n975), .Y(n1071) );
  INVX1_LVT U1231 ( .A(n1071), .Y(n1076) );
  AO22X1_LVT U1233 ( .A1(\regs[23][2] ), .A2(n968), .A3(\regs[12][2] ), .A4(
        n983), .Y(n1073) );
  INVX1_LVT U1234 ( .A(n1073), .Y(n1075) );
  NAND2X0_LVT U1235 ( .A1(\regs[29][2] ), .A2(n973), .Y(n1074) );
  NAND3X0_LVT U1236 ( .A1(n1076), .A2(n1075), .A3(n1074), .Y(n1105) );
  AO22X1_LVT U1239 ( .A1(\regs[16][2] ), .A2(n1003), .A3(\regs[20][2] ), .A4(
        n1001), .Y(n1084) );
  AO22X1_LVT U1241 ( .A1(\regs[27][2] ), .A2(n982), .A3(\regs[17][2] ), .A4(
        n990), .Y(n1083) );
  AO22X1_LVT U1243 ( .A1(\regs[10][2] ), .A2(n972), .A3(\regs[21][2] ), .A4(
        n969), .Y(n1082) );
  AO22X1_LVT U1245 ( .A1(\regs[15][2] ), .A2(n1015), .A3(\regs[24][2] ), .A4(
        n1005), .Y(n1081) );
  NOR4X1_LVT U1246 ( .A1(n1084), .A2(n1083), .A3(n1082), .A4(n1081), .Y(n1103)
         );
  AO22X1_LVT U1248 ( .A1(\regs[18][2] ), .A2(n995), .A3(\regs[13][2] ), .A4(
        n1025), .Y(n1092) );
  AO22X1_LVT U1250 ( .A1(\regs[3][2] ), .A2(n965), .A3(\regs[9][2] ), .A4(n967), .Y(n1091) );
  AO22X1_LVT U1252 ( .A1(\regs[14][2] ), .A2(n997), .A3(\regs[4][2] ), .A4(
        n1012), .Y(n1090) );
  AO22X1_LVT U1254 ( .A1(\regs[6][2] ), .A2(n1020), .A3(\regs[8][2] ), .A4(
        n981), .Y(n1089) );
  NOR4X1_LVT U1255 ( .A1(n1092), .A2(n1091), .A3(n1090), .A4(n1089), .Y(n1102)
         );
  AO22X1_LVT U1257 ( .A1(\regs[2][2] ), .A2(n1014), .A3(\regs[28][2] ), .A4(
        n986), .Y(n1100) );
  AO22X1_LVT U1258 ( .A1(\regs[31][2] ), .A2(n1027), .A3(\regs[25][2] ), .A4(
        n979), .Y(n1099) );
  AO22X1_LVT U1261 ( .A1(\regs[26][2] ), .A2(n1002), .A3(\regs[1][2] ), .A4(
        n998), .Y(n1098) );
  AO22X1_LVT U1263 ( .A1(\regs[11][2] ), .A2(n1022), .A3(\regs[19][2] ), .A4(
        n1017), .Y(n1097) );
  NOR4X1_LVT U1264 ( .A1(n1100), .A2(n1099), .A3(n1098), .A4(n1097), .Y(n1101)
         );
  NAND3X0_LVT U1265 ( .A1(n1103), .A2(n1102), .A3(n1101), .Y(n1104) );
  OR3X1_LVT U1266 ( .A1(n1106), .A2(n1105), .A3(n1104), .Y(n1107) );
  AO22X1_LVT U1267 ( .A1(wdata[2]), .A2(n960), .A3(n963), .A4(n1107), .Y(
        rdata1[2]) );
  AO22X1_LVT U1270 ( .A1(\regs[19][3] ), .A2(n1017), .A3(\regs[12][3] ), .A4(
        n983), .Y(n1144) );
  AO22X1_LVT U1272 ( .A1(\regs[22][3] ), .A2(n996), .A3(\regs[14][3] ), .A4(
        n997), .Y(n1112) );
  INVX1_LVT U1273 ( .A(n1112), .Y(n1117) );
  AO22X1_LVT U1275 ( .A1(\regs[2][3] ), .A2(n1014), .A3(\regs[7][3] ), .A4(
        n985), .Y(n1114) );
  INVX1_LVT U1276 ( .A(n1114), .Y(n1116) );
  NAND2X0_LVT U1277 ( .A1(\regs[11][3] ), .A2(n1022), .Y(n1115) );
  NAND3X0_LVT U1278 ( .A1(n1117), .A2(n1116), .A3(n1115), .Y(n1143) );
  AO22X1_LVT U1280 ( .A1(\regs[13][3] ), .A2(n1025), .A3(\regs[4][3] ), .A4(
        n1012), .Y(n1126) );
  AO22X1_LVT U1281 ( .A1(\regs[21][3] ), .A2(n969), .A3(\regs[6][3] ), .A4(
        n1020), .Y(n1125) );
  AO22X1_LVT U1283 ( .A1(\regs[31][3] ), .A2(n1027), .A3(\regs[18][3] ), .A4(
        n995), .Y(n1124) );
  AO22X1_LVT U1285 ( .A1(\regs[20][3] ), .A2(n1001), .A3(\regs[5][3] ), .A4(
        n987), .Y(n1123) );
  NOR4X1_LVT U1286 ( .A1(n1126), .A2(n1125), .A3(n1124), .A4(n1123), .Y(n1141)
         );
  AO22X1_LVT U1287 ( .A1(\regs[3][3] ), .A2(n965), .A3(\regs[1][3] ), .A4(n998), .Y(n1133) );
  AO22X1_LVT U1289 ( .A1(\regs[25][3] ), .A2(n979), .A3(\regs[28][3] ), .A4(
        n986), .Y(n1132) );
  AO22X1_LVT U1291 ( .A1(\regs[23][3] ), .A2(n968), .A3(\regs[17][3] ), .A4(
        n990), .Y(n1131) );
  AO22X1_LVT U1292 ( .A1(\regs[16][3] ), .A2(n1003), .A3(\regs[8][3] ), .A4(
        n981), .Y(n1130) );
  NOR4X1_LVT U1293 ( .A1(n1133), .A2(n1132), .A3(n1131), .A4(n1130), .Y(n1140)
         );
  AO22X1_LVT U1294 ( .A1(\regs[15][3] ), .A2(n1015), .A3(\regs[26][3] ), .A4(
        n1002), .Y(n1138) );
  AO22X1_LVT U1295 ( .A1(\regs[29][3] ), .A2(n973), .A3(\regs[24][3] ), .A4(
        n1005), .Y(n1137) );
  AO22X1_LVT U1296 ( .A1(\regs[27][3] ), .A2(n982), .A3(\regs[9][3] ), .A4(
        n967), .Y(n1136) );
  AO22X1_LVT U1297 ( .A1(\regs[30][3] ), .A2(n975), .A3(\regs[10][3] ), .A4(
        n972), .Y(n1135) );
  NOR4X1_LVT U1298 ( .A1(n1138), .A2(n1137), .A3(n1136), .A4(n1135), .Y(n1139)
         );
  NAND3X0_LVT U1299 ( .A1(n1141), .A2(n1140), .A3(n1139), .Y(n1142) );
  OR3X1_LVT U1300 ( .A1(n1144), .A2(n1143), .A3(n1142), .Y(n1145) );
  AO22X1_LVT U1301 ( .A1(wdata[3]), .A2(n960), .A3(n963), .A4(n1145), .Y(
        rdata1[3]) );
  AO22X1_LVT U1303 ( .A1(\regs[2][4] ), .A2(n1014), .A3(\regs[31][4] ), .A4(
        n1027), .Y(n1171) );
  AO22X1_LVT U1305 ( .A1(\regs[28][4] ), .A2(n986), .A3(\regs[16][4] ), .A4(
        n1003), .Y(n1146) );
  INVX1_LVT U1306 ( .A(n1146), .Y(n1151) );
  AO22X1_LVT U1307 ( .A1(\regs[13][4] ), .A2(n1025), .A3(\regs[25][4] ), .A4(
        n979), .Y(n1147) );
  INVX1_LVT U1308 ( .A(n1147), .Y(n1150) );
  NAND2X0_LVT U1310 ( .A1(\regs[15][4] ), .A2(n1015), .Y(n1149) );
  NAND3X0_LVT U1311 ( .A1(n1151), .A2(n1150), .A3(n1149), .Y(n1170) );
  AO22X1_LVT U1312 ( .A1(\regs[7][4] ), .A2(n985), .A3(\regs[30][4] ), .A4(
        n975), .Y(n1155) );
  AO22X1_LVT U1314 ( .A1(\regs[8][4] ), .A2(n981), .A3(\regs[29][4] ), .A4(
        n973), .Y(n1154) );
  AO22X1_LVT U1315 ( .A1(\regs[12][4] ), .A2(n983), .A3(\regs[9][4] ), .A4(
        n967), .Y(n1153) );
  AO22X1_LVT U1316 ( .A1(\regs[27][4] ), .A2(n982), .A3(\regs[18][4] ), .A4(
        n995), .Y(n1152) );
  NOR4X1_LVT U1317 ( .A1(n1155), .A2(n1154), .A3(n1153), .A4(n1152), .Y(n1168)
         );
  AO22X1_LVT U1318 ( .A1(\regs[26][4] ), .A2(n1002), .A3(\regs[17][4] ), .A4(
        n990), .Y(n1160) );
  AO22X1_LVT U1319 ( .A1(\regs[6][4] ), .A2(n1020), .A3(\regs[4][4] ), .A4(
        n1012), .Y(n1159) );
  AO22X1_LVT U1320 ( .A1(\regs[3][4] ), .A2(n965), .A3(\regs[24][4] ), .A4(
        n1005), .Y(n1158) );
  AO22X1_LVT U1321 ( .A1(\regs[23][4] ), .A2(n968), .A3(\regs[14][4] ), .A4(
        n997), .Y(n1157) );
  NOR4X1_LVT U1322 ( .A1(n1160), .A2(n1159), .A3(n1158), .A4(n1157), .Y(n1167)
         );
  AO22X1_LVT U1323 ( .A1(\regs[10][4] ), .A2(n972), .A3(\regs[19][4] ), .A4(
        n1017), .Y(n1165) );
  AO22X1_LVT U1324 ( .A1(\regs[20][4] ), .A2(n1001), .A3(\regs[5][4] ), .A4(
        n987), .Y(n1164) );
  AO22X1_LVT U1325 ( .A1(\regs[21][4] ), .A2(n969), .A3(\regs[1][4] ), .A4(
        n998), .Y(n1163) );
  AO22X1_LVT U1327 ( .A1(\regs[11][4] ), .A2(n1022), .A3(\regs[22][4] ), .A4(
        n996), .Y(n1162) );
  NOR4X1_LVT U1328 ( .A1(n1165), .A2(n1164), .A3(n1163), .A4(n1162), .Y(n1166)
         );
  NAND3X0_LVT U1329 ( .A1(n1168), .A2(n1167), .A3(n1166), .Y(n1169) );
  OR3X1_LVT U1330 ( .A1(n1171), .A2(n1170), .A3(n1169), .Y(n1172) );
  AO22X1_LVT U1331 ( .A1(wdata[4]), .A2(n960), .A3(n963), .A4(n1172), .Y(
        rdata1[4]) );
  AO22X1_LVT U1333 ( .A1(\regs[5][5] ), .A2(n987), .A3(\regs[9][5] ), .A4(n967), .Y(n1197) );
  AO22X1_LVT U1334 ( .A1(\regs[7][5] ), .A2(n985), .A3(\regs[29][5] ), .A4(
        n973), .Y(n1173) );
  INVX1_LVT U1335 ( .A(n1173), .Y(n1177) );
  AO22X1_LVT U1336 ( .A1(\regs[23][5] ), .A2(n968), .A3(\regs[14][5] ), .A4(
        n997), .Y(n1174) );
  INVX1_LVT U1337 ( .A(n1174), .Y(n1176) );
  NAND2X0_LVT U1338 ( .A1(\regs[31][5] ), .A2(n1027), .Y(n1175) );
  NAND3X0_LVT U1339 ( .A1(n1177), .A2(n1176), .A3(n1175), .Y(n1196) );
  AO22X1_LVT U1340 ( .A1(\regs[12][5] ), .A2(n983), .A3(\regs[21][5] ), .A4(
        n969), .Y(n1181) );
  AO22X1_LVT U1341 ( .A1(\regs[19][5] ), .A2(n1017), .A3(\regs[2][5] ), .A4(
        n1014), .Y(n1180) );
  AO22X1_LVT U1342 ( .A1(\regs[25][5] ), .A2(n979), .A3(\regs[8][5] ), .A4(
        n981), .Y(n1179) );
  AO22X1_LVT U1343 ( .A1(\regs[20][5] ), .A2(n1001), .A3(\regs[17][5] ), .A4(
        n990), .Y(n1178) );
  NOR4X1_LVT U1344 ( .A1(n1181), .A2(n1180), .A3(n1179), .A4(n1178), .Y(n1194)
         );
  AO22X1_LVT U1345 ( .A1(\regs[10][5] ), .A2(n972), .A3(\regs[4][5] ), .A4(
        n1012), .Y(n1185) );
  AO22X1_LVT U1346 ( .A1(\regs[30][5] ), .A2(n975), .A3(\regs[6][5] ), .A4(
        n1020), .Y(n1184) );
  AO22X1_LVT U1347 ( .A1(\regs[27][5] ), .A2(n982), .A3(\regs[1][5] ), .A4(
        n998), .Y(n1183) );
  AO22X1_LVT U1348 ( .A1(\regs[3][5] ), .A2(n965), .A3(\regs[11][5] ), .A4(
        n1022), .Y(n1182) );
  NOR4X1_LVT U1349 ( .A1(n1185), .A2(n1184), .A3(n1183), .A4(n1182), .Y(n1193)
         );
  AO22X1_LVT U1350 ( .A1(\regs[26][5] ), .A2(n1002), .A3(\regs[18][5] ), .A4(
        n995), .Y(n1191) );
  AO22X1_LVT U1352 ( .A1(\regs[28][5] ), .A2(n986), .A3(\regs[22][5] ), .A4(
        n996), .Y(n1190) );
  AO22X1_LVT U1353 ( .A1(\regs[13][5] ), .A2(n1025), .A3(\regs[24][5] ), .A4(
        n1005), .Y(n1189) );
  AO22X1_LVT U1354 ( .A1(\regs[15][5] ), .A2(n1015), .A3(\regs[16][5] ), .A4(
        n1003), .Y(n1188) );
  NOR4X1_LVT U1355 ( .A1(n1191), .A2(n1190), .A3(n1189), .A4(n1188), .Y(n1192)
         );
  NAND3X0_LVT U1356 ( .A1(n1194), .A2(n1193), .A3(n1192), .Y(n1195) );
  OR3X1_LVT U1357 ( .A1(n1197), .A2(n1196), .A3(n1195), .Y(n1198) );
  AO22X1_LVT U1358 ( .A1(wdata[5]), .A2(n960), .A3(n963), .A4(n1198), .Y(
        rdata1[5]) );
  AO22X1_LVT U1360 ( .A1(\regs[15][6] ), .A2(n1015), .A3(\regs[22][6] ), .A4(
        n996), .Y(n1224) );
  AO22X1_LVT U1361 ( .A1(\regs[30][6] ), .A2(n975), .A3(\regs[26][6] ), .A4(
        n1002), .Y(n1199) );
  INVX1_LVT U1362 ( .A(n1199), .Y(n1204) );
  AO22X1_LVT U1364 ( .A1(\regs[4][6] ), .A2(n1012), .A3(\regs[24][6] ), .A4(
        n1005), .Y(n1201) );
  INVX1_LVT U1365 ( .A(n1201), .Y(n1203) );
  NAND2X0_LVT U1366 ( .A1(\regs[16][6] ), .A2(n1003), .Y(n1202) );
  NAND3X0_LVT U1367 ( .A1(n1204), .A2(n1203), .A3(n1202), .Y(n1223) );
  AO22X1_LVT U1368 ( .A1(\regs[12][6] ), .A2(n983), .A3(\regs[6][6] ), .A4(
        n1020), .Y(n1208) );
  AO22X1_LVT U1369 ( .A1(\regs[2][6] ), .A2(n1014), .A3(\regs[21][6] ), .A4(
        n969), .Y(n1207) );
  AO22X1_LVT U1370 ( .A1(\regs[19][6] ), .A2(n1017), .A3(\regs[17][6] ), .A4(
        n990), .Y(n1206) );
  AO22X1_LVT U1371 ( .A1(\regs[7][6] ), .A2(n985), .A3(\regs[18][6] ), .A4(
        n995), .Y(n1205) );
  NOR4X1_LVT U1372 ( .A1(n1208), .A2(n1207), .A3(n1206), .A4(n1205), .Y(n1221)
         );
  AO22X1_LVT U1373 ( .A1(\regs[13][6] ), .A2(n1025), .A3(\regs[3][6] ), .A4(
        n965), .Y(n1213) );
  AO22X1_LVT U1375 ( .A1(\regs[8][6] ), .A2(n981), .A3(\regs[25][6] ), .A4(
        n979), .Y(n1212) );
  AO22X1_LVT U1376 ( .A1(\regs[5][6] ), .A2(n987), .A3(\regs[9][6] ), .A4(n967), .Y(n1211) );
  AO22X1_LVT U1377 ( .A1(\regs[14][6] ), .A2(n997), .A3(\regs[28][6] ), .A4(
        n986), .Y(n1210) );
  NOR4X1_LVT U1378 ( .A1(n1213), .A2(n1212), .A3(n1211), .A4(n1210), .Y(n1220)
         );
  AO22X1_LVT U1379 ( .A1(\regs[10][6] ), .A2(n972), .A3(\regs[23][6] ), .A4(
        n968), .Y(n1218) );
  AO22X1_LVT U1381 ( .A1(\regs[29][6] ), .A2(n973), .A3(\regs[27][6] ), .A4(
        n982), .Y(n1217) );
  AO22X1_LVT U1382 ( .A1(\regs[11][6] ), .A2(n1022), .A3(\regs[31][6] ), .A4(
        n1027), .Y(n1216) );
  AO22X1_LVT U1383 ( .A1(\regs[20][6] ), .A2(n1001), .A3(\regs[1][6] ), .A4(
        n998), .Y(n1215) );
  NOR4X1_LVT U1384 ( .A1(n1218), .A2(n1217), .A3(n1216), .A4(n1215), .Y(n1219)
         );
  NAND3X0_LVT U1385 ( .A1(n1221), .A2(n1220), .A3(n1219), .Y(n1222) );
  OR3X1_LVT U1386 ( .A1(n1224), .A2(n1223), .A3(n1222), .Y(n1225) );
  AO22X1_LVT U1387 ( .A1(wdata[6]), .A2(n960), .A3(n963), .A4(n1225), .Y(
        rdata1[6]) );
  AO22X1_LVT U1389 ( .A1(\regs[19][7] ), .A2(n1017), .A3(\regs[30][7] ), .A4(
        n975), .Y(n1250) );
  AO22X1_LVT U1390 ( .A1(\regs[4][7] ), .A2(n1012), .A3(\regs[3][7] ), .A4(
        n965), .Y(n1227) );
  INVX1_LVT U1391 ( .A(n1227), .Y(n1231) );
  AO22X1_LVT U1392 ( .A1(\regs[2][7] ), .A2(n1014), .A3(\regs[10][7] ), .A4(
        n972), .Y(n1228) );
  INVX1_LVT U1393 ( .A(n1228), .Y(n1230) );
  NAND2X0_LVT U1394 ( .A1(\regs[12][7] ), .A2(n983), .Y(n1229) );
  NAND3X0_LVT U1395 ( .A1(n1231), .A2(n1230), .A3(n1229), .Y(n1249) );
  AO22X1_LVT U1396 ( .A1(\regs[11][7] ), .A2(n1022), .A3(\regs[14][7] ), .A4(
        n997), .Y(n1235) );
  AO22X1_LVT U1397 ( .A1(\regs[18][7] ), .A2(n995), .A3(\regs[27][7] ), .A4(
        n982), .Y(n1234) );
  AO22X1_LVT U1398 ( .A1(\regs[28][7] ), .A2(n986), .A3(\regs[17][7] ), .A4(
        n990), .Y(n1233) );
  AO22X1_LVT U1399 ( .A1(\regs[16][7] ), .A2(n1003), .A3(\regs[9][7] ), .A4(
        n967), .Y(n1232) );
  NOR4X1_LVT U1400 ( .A1(n1235), .A2(n1234), .A3(n1233), .A4(n1232), .Y(n1247)
         );
  AO22X1_LVT U1401 ( .A1(\regs[8][7] ), .A2(n981), .A3(\regs[22][7] ), .A4(
        n996), .Y(n1240) );
  AO22X1_LVT U1402 ( .A1(\regs[23][7] ), .A2(n968), .A3(\regs[21][7] ), .A4(
        n969), .Y(n1239) );
  AO22X1_LVT U1403 ( .A1(\regs[24][7] ), .A2(n1005), .A3(\regs[5][7] ), .A4(
        n987), .Y(n1238) );
  AO22X1_LVT U1404 ( .A1(\regs[29][7] ), .A2(n973), .A3(\regs[25][7] ), .A4(
        n979), .Y(n1237) );
  NOR4X1_LVT U1405 ( .A1(n1240), .A2(n1239), .A3(n1238), .A4(n1237), .Y(n1246)
         );
  AO22X1_LVT U1406 ( .A1(\regs[1][7] ), .A2(n998), .A3(\regs[15][7] ), .A4(
        n1015), .Y(n1244) );
  AO22X1_LVT U1407 ( .A1(\regs[20][7] ), .A2(n1001), .A3(\regs[13][7] ), .A4(
        n1025), .Y(n1243) );
  AO22X1_LVT U1408 ( .A1(\regs[6][7] ), .A2(n1020), .A3(\regs[31][7] ), .A4(
        n1027), .Y(n1242) );
  AO22X1_LVT U1409 ( .A1(\regs[26][7] ), .A2(n1002), .A3(\regs[7][7] ), .A4(
        n985), .Y(n1241) );
  NOR4X1_LVT U1410 ( .A1(n1244), .A2(n1243), .A3(n1242), .A4(n1241), .Y(n1245)
         );
  NAND3X0_LVT U1411 ( .A1(n1247), .A2(n1246), .A3(n1245), .Y(n1248) );
  OR3X1_LVT U1412 ( .A1(n1250), .A2(n1249), .A3(n1248), .Y(n1251) );
  AO22X1_LVT U1413 ( .A1(wdata[7]), .A2(n960), .A3(n963), .A4(n1251), .Y(
        rdata1[7]) );
  AO22X1_LVT U1415 ( .A1(\regs[20][8] ), .A2(n1001), .A3(\regs[14][8] ), .A4(
        n997), .Y(n1275) );
  AO22X1_LVT U1416 ( .A1(\regs[8][8] ), .A2(n981), .A3(\regs[6][8] ), .A4(
        n1020), .Y(n1252) );
  INVX1_LVT U1417 ( .A(n1252), .Y(n1256) );
  AO22X1_LVT U1418 ( .A1(\regs[28][8] ), .A2(n986), .A3(\regs[7][8] ), .A4(
        n985), .Y(n1253) );
  INVX1_LVT U1419 ( .A(n1253), .Y(n1255) );
  NAND2X0_LVT U1420 ( .A1(\regs[12][8] ), .A2(n983), .Y(n1254) );
  NAND3X0_LVT U1421 ( .A1(n1256), .A2(n1255), .A3(n1254), .Y(n1274) );
  AO22X1_LVT U1422 ( .A1(\regs[31][8] ), .A2(n1027), .A3(\regs[13][8] ), .A4(
        n1025), .Y(n1260) );
  AO22X1_LVT U1423 ( .A1(\regs[23][8] ), .A2(n968), .A3(\regs[30][8] ), .A4(
        n975), .Y(n1259) );
  AO22X1_LVT U1424 ( .A1(\regs[5][8] ), .A2(n987), .A3(\regs[16][8] ), .A4(
        n1003), .Y(n1258) );
  AO22X1_LVT U1425 ( .A1(\regs[15][8] ), .A2(n1015), .A3(\regs[4][8] ), .A4(
        n1012), .Y(n1257) );
  NOR4X1_LVT U1426 ( .A1(n1260), .A2(n1259), .A3(n1258), .A4(n1257), .Y(n1272)
         );
  AO22X1_LVT U1427 ( .A1(\regs[27][8] ), .A2(n982), .A3(\regs[29][8] ), .A4(
        n973), .Y(n1264) );
  AO22X1_LVT U1428 ( .A1(\regs[22][8] ), .A2(n996), .A3(\regs[1][8] ), .A4(
        n998), .Y(n1263) );
  AO22X1_LVT U1429 ( .A1(\regs[18][8] ), .A2(n995), .A3(\regs[17][8] ), .A4(
        n990), .Y(n1262) );
  AO22X1_LVT U1430 ( .A1(\regs[10][8] ), .A2(n972), .A3(\regs[25][8] ), .A4(
        n979), .Y(n1261) );
  NOR4X1_LVT U1431 ( .A1(n1264), .A2(n1263), .A3(n1262), .A4(n1261), .Y(n1271)
         );
  AO22X1_LVT U1432 ( .A1(\regs[24][8] ), .A2(n1005), .A3(\regs[26][8] ), .A4(
        n1002), .Y(n1269) );
  AO22X1_LVT U1433 ( .A1(\regs[19][8] ), .A2(n1017), .A3(\regs[2][8] ), .A4(
        n1014), .Y(n1268) );
  AO22X1_LVT U1435 ( .A1(\regs[9][8] ), .A2(n967), .A3(\regs[3][8] ), .A4(n965), .Y(n1267) );
  AO22X1_LVT U1436 ( .A1(\regs[11][8] ), .A2(n1022), .A3(\regs[21][8] ), .A4(
        n969), .Y(n1266) );
  NOR4X1_LVT U1437 ( .A1(n1269), .A2(n1268), .A3(n1267), .A4(n1266), .Y(n1270)
         );
  NAND3X0_LVT U1438 ( .A1(n1272), .A2(n1271), .A3(n1270), .Y(n1273) );
  OR3X1_LVT U1439 ( .A1(n1275), .A2(n1274), .A3(n1273), .Y(n1276) );
  AO22X1_LVT U1440 ( .A1(wdata[8]), .A2(n960), .A3(n963), .A4(n1276), .Y(
        rdata1[8]) );
  AO22X1_LVT U1442 ( .A1(\regs[23][9] ), .A2(n968), .A3(\regs[24][9] ), .A4(
        n1005), .Y(n1299) );
  AO22X1_LVT U1443 ( .A1(\regs[15][9] ), .A2(n1015), .A3(\regs[8][9] ), .A4(
        n981), .Y(n1277) );
  INVX1_LVT U1444 ( .A(n1277), .Y(n1281) );
  AO22X1_LVT U1445 ( .A1(\regs[26][9] ), .A2(n1002), .A3(\regs[29][9] ), .A4(
        n973), .Y(n1278) );
  INVX1_LVT U1446 ( .A(n1278), .Y(n1280) );
  NAND2X0_LVT U1447 ( .A1(\regs[1][9] ), .A2(n998), .Y(n1279) );
  NAND3X0_LVT U1448 ( .A1(n1281), .A2(n1280), .A3(n1279), .Y(n1298) );
  AO22X1_LVT U1449 ( .A1(\regs[12][9] ), .A2(n983), .A3(\regs[16][9] ), .A4(
        n1003), .Y(n1285) );
  AO22X1_LVT U1450 ( .A1(\regs[9][9] ), .A2(n967), .A3(\regs[17][9] ), .A4(
        n990), .Y(n1284) );
  AO22X1_LVT U1451 ( .A1(\regs[28][9] ), .A2(n986), .A3(\regs[2][9] ), .A4(
        n1014), .Y(n1283) );
  AO22X1_LVT U1452 ( .A1(\regs[14][9] ), .A2(n997), .A3(\regs[7][9] ), .A4(
        n985), .Y(n1282) );
  NOR4X1_LVT U1453 ( .A1(n1285), .A2(n1284), .A3(n1283), .A4(n1282), .Y(n1296)
         );
  AO22X1_LVT U1454 ( .A1(\regs[6][9] ), .A2(n1020), .A3(\regs[31][9] ), .A4(
        n1027), .Y(n1289) );
  AO22X1_LVT U1455 ( .A1(\regs[21][9] ), .A2(n969), .A3(\regs[4][9] ), .A4(
        n1012), .Y(n1288) );
  AO22X1_LVT U1456 ( .A1(\regs[5][9] ), .A2(n987), .A3(\regs[30][9] ), .A4(
        n975), .Y(n1287) );
  AO22X1_LVT U1457 ( .A1(\regs[27][9] ), .A2(n982), .A3(\regs[19][9] ), .A4(
        n1017), .Y(n1286) );
  NOR4X1_LVT U1458 ( .A1(n1289), .A2(n1288), .A3(n1287), .A4(n1286), .Y(n1295)
         );
  AO22X1_LVT U1459 ( .A1(\regs[11][9] ), .A2(n1022), .A3(\regs[3][9] ), .A4(
        n965), .Y(n1293) );
  AO22X1_LVT U1460 ( .A1(\regs[20][9] ), .A2(n1001), .A3(\regs[18][9] ), .A4(
        n995), .Y(n1292) );
  AO22X1_LVT U1461 ( .A1(\regs[22][9] ), .A2(n996), .A3(\regs[13][9] ), .A4(
        n1025), .Y(n1291) );
  AO22X1_LVT U1462 ( .A1(\regs[25][9] ), .A2(n979), .A3(\regs[10][9] ), .A4(
        n972), .Y(n1290) );
  NOR4X1_LVT U1463 ( .A1(n1293), .A2(n1292), .A3(n1291), .A4(n1290), .Y(n1294)
         );
  NAND3X0_LVT U1464 ( .A1(n1296), .A2(n1295), .A3(n1294), .Y(n1297) );
  OR3X1_LVT U1465 ( .A1(n1299), .A2(n1298), .A3(n1297), .Y(n1300) );
  AO22X1_LVT U1466 ( .A1(wdata[9]), .A2(n960), .A3(n963), .A4(n1300), .Y(
        rdata1[9]) );
  AO22X1_LVT U1468 ( .A1(\regs[8][10] ), .A2(n981), .A3(\regs[26][10] ), .A4(
        n1002), .Y(n1323) );
  AO22X1_LVT U1469 ( .A1(\regs[22][10] ), .A2(n996), .A3(\regs[18][10] ), .A4(
        n995), .Y(n1301) );
  INVX1_LVT U1470 ( .A(n1301), .Y(n1305) );
  AO22X1_LVT U1471 ( .A1(\regs[17][10] ), .A2(n990), .A3(\regs[11][10] ), .A4(
        n1022), .Y(n1302) );
  INVX1_LVT U1472 ( .A(n1302), .Y(n1304) );
  NAND2X0_LVT U1473 ( .A1(\regs[2][10] ), .A2(n1014), .Y(n1303) );
  NAND3X0_LVT U1474 ( .A1(n1305), .A2(n1304), .A3(n1303), .Y(n1322) );
  AO22X1_LVT U1475 ( .A1(\regs[24][10] ), .A2(n1005), .A3(\regs[13][10] ), 
        .A4(n1025), .Y(n1309) );
  AO22X1_LVT U1476 ( .A1(\regs[9][10] ), .A2(n967), .A3(\regs[27][10] ), .A4(
        n982), .Y(n1308) );
  AO22X1_LVT U1477 ( .A1(\regs[5][10] ), .A2(n987), .A3(\regs[31][10] ), .A4(
        n1027), .Y(n1307) );
  AO22X1_LVT U1478 ( .A1(\regs[30][10] ), .A2(n975), .A3(\regs[16][10] ), .A4(
        n1003), .Y(n1306) );
  NOR4X1_LVT U1479 ( .A1(n1309), .A2(n1308), .A3(n1307), .A4(n1306), .Y(n1320)
         );
  AO22X1_LVT U1480 ( .A1(\regs[12][10] ), .A2(n983), .A3(\regs[28][10] ), .A4(
        n986), .Y(n1313) );
  AO22X1_LVT U1481 ( .A1(\regs[3][10] ), .A2(n965), .A3(\regs[19][10] ), .A4(
        n1017), .Y(n1312) );
  AO22X1_LVT U1482 ( .A1(\regs[6][10] ), .A2(n1020), .A3(\regs[15][10] ), .A4(
        n1015), .Y(n1311) );
  AO22X1_LVT U1483 ( .A1(\regs[21][10] ), .A2(n969), .A3(\regs[20][10] ), .A4(
        n1001), .Y(n1310) );
  NOR4X1_LVT U1484 ( .A1(n1313), .A2(n1312), .A3(n1311), .A4(n1310), .Y(n1319)
         );
  AO22X1_LVT U1485 ( .A1(\regs[29][10] ), .A2(n973), .A3(\regs[23][10] ), .A4(
        n968), .Y(n1317) );
  AO22X1_LVT U1486 ( .A1(\regs[7][10] ), .A2(n985), .A3(\regs[4][10] ), .A4(
        n1012), .Y(n1316) );
  AO22X1_LVT U1487 ( .A1(\regs[14][10] ), .A2(n997), .A3(\regs[10][10] ), .A4(
        n972), .Y(n1315) );
  AO22X1_LVT U1488 ( .A1(\regs[1][10] ), .A2(n998), .A3(\regs[25][10] ), .A4(
        n979), .Y(n1314) );
  NOR4X1_LVT U1489 ( .A1(n1317), .A2(n1316), .A3(n1315), .A4(n1314), .Y(n1318)
         );
  NAND3X0_LVT U1490 ( .A1(n1320), .A2(n1319), .A3(n1318), .Y(n1321) );
  OR3X1_LVT U1491 ( .A1(n1323), .A2(n1322), .A3(n1321), .Y(n1324) );
  AO22X1_LVT U1492 ( .A1(wdata[10]), .A2(n960), .A3(n963), .A4(n1324), .Y(
        rdata1[10]) );
  AO22X1_LVT U1495 ( .A1(\regs[22][11] ), .A2(n996), .A3(\regs[7][11] ), .A4(
        n985), .Y(n1348) );
  AO22X1_LVT U1496 ( .A1(\regs[27][11] ), .A2(n982), .A3(\regs[21][11] ), .A4(
        n969), .Y(n1326) );
  INVX1_LVT U1497 ( .A(n1326), .Y(n1330) );
  AO22X1_LVT U1498 ( .A1(\regs[30][11] ), .A2(n975), .A3(\regs[20][11] ), .A4(
        n1001), .Y(n1327) );
  INVX1_LVT U1499 ( .A(n1327), .Y(n1329) );
  NAND2X0_LVT U1500 ( .A1(\regs[18][11] ), .A2(n995), .Y(n1328) );
  NAND3X0_LVT U1501 ( .A1(n1330), .A2(n1329), .A3(n1328), .Y(n1347) );
  AO22X1_LVT U1502 ( .A1(\regs[19][11] ), .A2(n1017), .A3(\regs[9][11] ), .A4(
        n967), .Y(n1334) );
  AO22X1_LVT U1503 ( .A1(\regs[2][11] ), .A2(n1014), .A3(\regs[3][11] ), .A4(
        n965), .Y(n1333) );
  AO22X1_LVT U1504 ( .A1(\regs[6][11] ), .A2(n1020), .A3(\regs[31][11] ), .A4(
        n1027), .Y(n1332) );
  AO22X1_LVT U1505 ( .A1(\regs[5][11] ), .A2(n987), .A3(\regs[1][11] ), .A4(
        n998), .Y(n1331) );
  NOR4X1_LVT U1506 ( .A1(n1334), .A2(n1333), .A3(n1332), .A4(n1331), .Y(n1345)
         );
  AO22X1_LVT U1507 ( .A1(\regs[13][11] ), .A2(n1025), .A3(\regs[12][11] ), 
        .A4(n983), .Y(n1338) );
  AO22X1_LVT U1508 ( .A1(\regs[15][11] ), .A2(n1015), .A3(\regs[11][11] ), 
        .A4(n1022), .Y(n1337) );
  AO22X1_LVT U1509 ( .A1(\regs[25][11] ), .A2(n979), .A3(\regs[23][11] ), .A4(
        n968), .Y(n1336) );
  AO22X1_LVT U1510 ( .A1(\regs[8][11] ), .A2(n981), .A3(\regs[4][11] ), .A4(
        n1012), .Y(n1335) );
  NOR4X1_LVT U1511 ( .A1(n1338), .A2(n1337), .A3(n1336), .A4(n1335), .Y(n1344)
         );
  AO22X1_LVT U1512 ( .A1(\regs[10][11] ), .A2(n972), .A3(\regs[29][11] ), .A4(
        n973), .Y(n1342) );
  AO22X1_LVT U1513 ( .A1(\regs[28][11] ), .A2(n986), .A3(\regs[17][11] ), .A4(
        n990), .Y(n1341) );
  AO22X1_LVT U1514 ( .A1(\regs[26][11] ), .A2(n1002), .A3(\regs[14][11] ), 
        .A4(n997), .Y(n1340) );
  AO22X1_LVT U1515 ( .A1(\regs[24][11] ), .A2(n1005), .A3(\regs[16][11] ), 
        .A4(n1003), .Y(n1339) );
  NOR4X1_LVT U1516 ( .A1(n1342), .A2(n1341), .A3(n1340), .A4(n1339), .Y(n1343)
         );
  NAND3X0_LVT U1517 ( .A1(n1345), .A2(n1344), .A3(n1343), .Y(n1346) );
  OR3X1_LVT U1518 ( .A1(n1348), .A2(n1347), .A3(n1346), .Y(n1349) );
  AO22X1_LVT U1519 ( .A1(wdata[11]), .A2(n960), .A3(n963), .A4(n1349), .Y(
        rdata1[11]) );
  AO22X1_LVT U1521 ( .A1(\regs[31][12] ), .A2(n1027), .A3(\regs[5][12] ), .A4(
        n987), .Y(n1372) );
  AO22X1_LVT U1522 ( .A1(\regs[2][12] ), .A2(n1014), .A3(\regs[4][12] ), .A4(
        n1012), .Y(n1350) );
  INVX1_LVT U1523 ( .A(n1350), .Y(n1354) );
  AO22X1_LVT U1524 ( .A1(\regs[19][12] ), .A2(n1017), .A3(\regs[18][12] ), 
        .A4(n995), .Y(n1351) );
  INVX1_LVT U1525 ( .A(n1351), .Y(n1353) );
  NAND2X0_LVT U1526 ( .A1(\regs[29][12] ), .A2(n973), .Y(n1352) );
  NAND3X0_LVT U1527 ( .A1(n1354), .A2(n1353), .A3(n1352), .Y(n1371) );
  AO22X1_LVT U1528 ( .A1(\regs[21][12] ), .A2(n969), .A3(\regs[28][12] ), .A4(
        n986), .Y(n1358) );
  AO22X1_LVT U1529 ( .A1(\regs[24][12] ), .A2(n1005), .A3(\regs[23][12] ), 
        .A4(n968), .Y(n1357) );
  AO22X1_LVT U1530 ( .A1(\regs[22][12] ), .A2(n996), .A3(\regs[30][12] ), .A4(
        n975), .Y(n1356) );
  AO22X1_LVT U1531 ( .A1(\regs[16][12] ), .A2(n1003), .A3(\regs[6][12] ), .A4(
        n1020), .Y(n1355) );
  NOR4X1_LVT U1532 ( .A1(n1358), .A2(n1357), .A3(n1356), .A4(n1355), .Y(n1369)
         );
  AO22X1_LVT U1533 ( .A1(\regs[20][12] ), .A2(n1001), .A3(\regs[26][12] ), 
        .A4(n1002), .Y(n1362) );
  AO22X1_LVT U1534 ( .A1(\regs[15][12] ), .A2(n1015), .A3(\regs[9][12] ), .A4(
        n967), .Y(n1361) );
  AO22X1_LVT U1535 ( .A1(\regs[11][12] ), .A2(n1022), .A3(\regs[13][12] ), 
        .A4(n1025), .Y(n1360) );
  AO22X1_LVT U1536 ( .A1(\regs[12][12] ), .A2(n983), .A3(\regs[8][12] ), .A4(
        n981), .Y(n1359) );
  NOR4X1_LVT U1537 ( .A1(n1362), .A2(n1361), .A3(n1360), .A4(n1359), .Y(n1368)
         );
  AO22X1_LVT U1538 ( .A1(\regs[1][12] ), .A2(n998), .A3(\regs[17][12] ), .A4(
        n990), .Y(n1366) );
  AO22X1_LVT U1539 ( .A1(\regs[14][12] ), .A2(n997), .A3(\regs[10][12] ), .A4(
        n972), .Y(n1365) );
  AO22X1_LVT U1540 ( .A1(\regs[3][12] ), .A2(n965), .A3(\regs[27][12] ), .A4(
        n982), .Y(n1364) );
  AO22X1_LVT U1541 ( .A1(\regs[25][12] ), .A2(n979), .A3(\regs[7][12] ), .A4(
        n985), .Y(n1363) );
  NOR4X1_LVT U1542 ( .A1(n1366), .A2(n1365), .A3(n1364), .A4(n1363), .Y(n1367)
         );
  NAND3X0_LVT U1543 ( .A1(n1369), .A2(n1368), .A3(n1367), .Y(n1370) );
  OR3X1_LVT U1544 ( .A1(n1372), .A2(n1371), .A3(n1370), .Y(n1373) );
  AO22X1_LVT U1545 ( .A1(wdata[12]), .A2(n960), .A3(n963), .A4(n1373), .Y(
        rdata1[12]) );
  AO22X1_LVT U1547 ( .A1(\regs[29][13] ), .A2(n973), .A3(\regs[4][13] ), .A4(
        n1012), .Y(n1396) );
  AO22X1_LVT U1548 ( .A1(\regs[1][13] ), .A2(n998), .A3(\regs[11][13] ), .A4(
        n1022), .Y(n1374) );
  INVX1_LVT U1549 ( .A(n1374), .Y(n1378) );
  AO22X1_LVT U1550 ( .A1(\regs[15][13] ), .A2(n1015), .A3(\regs[20][13] ), 
        .A4(n1001), .Y(n1375) );
  INVX1_LVT U1551 ( .A(n1375), .Y(n1377) );
  NAND2X0_LVT U1552 ( .A1(\regs[9][13] ), .A2(n967), .Y(n1376) );
  NAND3X0_LVT U1553 ( .A1(n1378), .A2(n1377), .A3(n1376), .Y(n1395) );
  AO22X1_LVT U1554 ( .A1(\regs[25][13] ), .A2(n979), .A3(\regs[28][13] ), .A4(
        n986), .Y(n1382) );
  AO22X1_LVT U1555 ( .A1(\regs[14][13] ), .A2(n997), .A3(\regs[30][13] ), .A4(
        n975), .Y(n1381) );
  AO22X1_LVT U1556 ( .A1(\regs[12][13] ), .A2(n983), .A3(\regs[19][13] ), .A4(
        n1017), .Y(n1380) );
  AO22X1_LVT U1557 ( .A1(\regs[23][13] ), .A2(n968), .A3(\regs[18][13] ), .A4(
        n995), .Y(n1379) );
  NOR4X1_LVT U1558 ( .A1(n1382), .A2(n1381), .A3(n1380), .A4(n1379), .Y(n1393)
         );
  AO22X1_LVT U1559 ( .A1(\regs[16][13] ), .A2(n1003), .A3(\regs[27][13] ), 
        .A4(n982), .Y(n1386) );
  AO22X1_LVT U1560 ( .A1(\regs[8][13] ), .A2(n981), .A3(\regs[26][13] ), .A4(
        n1002), .Y(n1385) );
  AO22X1_LVT U1561 ( .A1(\regs[10][13] ), .A2(n972), .A3(\regs[7][13] ), .A4(
        n985), .Y(n1384) );
  AO22X1_LVT U1562 ( .A1(\regs[5][13] ), .A2(n987), .A3(\regs[21][13] ), .A4(
        n969), .Y(n1383) );
  NOR4X1_LVT U1563 ( .A1(n1386), .A2(n1385), .A3(n1384), .A4(n1383), .Y(n1392)
         );
  AO22X1_LVT U1564 ( .A1(\regs[24][13] ), .A2(n1005), .A3(\regs[13][13] ), 
        .A4(n1025), .Y(n1390) );
  AO22X1_LVT U1565 ( .A1(\regs[22][13] ), .A2(n996), .A3(\regs[3][13] ), .A4(
        n965), .Y(n1389) );
  AO22X1_LVT U1566 ( .A1(\regs[6][13] ), .A2(n1020), .A3(\regs[31][13] ), .A4(
        n1027), .Y(n1388) );
  AO22X1_LVT U1567 ( .A1(\regs[2][13] ), .A2(n1014), .A3(\regs[17][13] ), .A4(
        n990), .Y(n1387) );
  NOR4X1_LVT U1568 ( .A1(n1390), .A2(n1389), .A3(n1388), .A4(n1387), .Y(n1391)
         );
  NAND3X0_LVT U1569 ( .A1(n1393), .A2(n1392), .A3(n1391), .Y(n1394) );
  OR3X1_LVT U1570 ( .A1(n1396), .A2(n1395), .A3(n1394), .Y(n1397) );
  AO22X1_LVT U1571 ( .A1(wdata[13]), .A2(n960), .A3(n963), .A4(n1397), .Y(
        rdata1[13]) );
  AO22X1_LVT U1573 ( .A1(\regs[31][14] ), .A2(n1027), .A3(\regs[27][14] ), 
        .A4(n982), .Y(n1420) );
  AO22X1_LVT U1574 ( .A1(\regs[6][14] ), .A2(n1020), .A3(\regs[22][14] ), .A4(
        n996), .Y(n1398) );
  INVX1_LVT U1575 ( .A(n1398), .Y(n1402) );
  AO22X1_LVT U1576 ( .A1(\regs[15][14] ), .A2(n1015), .A3(\regs[2][14] ), .A4(
        n1014), .Y(n1399) );
  INVX1_LVT U1577 ( .A(n1399), .Y(n1401) );
  NAND2X0_LVT U1578 ( .A1(\regs[23][14] ), .A2(n968), .Y(n1400) );
  NAND3X0_LVT U1579 ( .A1(n1402), .A2(n1401), .A3(n1400), .Y(n1419) );
  AO22X1_LVT U1580 ( .A1(\regs[19][14] ), .A2(n1017), .A3(\regs[10][14] ), 
        .A4(n972), .Y(n1406) );
  AO22X1_LVT U1581 ( .A1(\regs[3][14] ), .A2(n965), .A3(\regs[4][14] ), .A4(
        n1012), .Y(n1405) );
  AO22X1_LVT U1582 ( .A1(\regs[8][14] ), .A2(n981), .A3(\regs[7][14] ), .A4(
        n985), .Y(n1404) );
  AO22X1_LVT U1583 ( .A1(\regs[28][14] ), .A2(n986), .A3(\regs[12][14] ), .A4(
        n983), .Y(n1403) );
  NOR4X1_LVT U1584 ( .A1(n1406), .A2(n1405), .A3(n1404), .A4(n1403), .Y(n1417)
         );
  AO22X1_LVT U1585 ( .A1(\regs[25][14] ), .A2(n979), .A3(\regs[21][14] ), .A4(
        n969), .Y(n1410) );
  AO22X1_LVT U1586 ( .A1(\regs[18][14] ), .A2(n995), .A3(\regs[9][14] ), .A4(
        n967), .Y(n1409) );
  AO22X1_LVT U1587 ( .A1(\regs[24][14] ), .A2(n1005), .A3(\regs[14][14] ), 
        .A4(n997), .Y(n1408) );
  AO22X1_LVT U1588 ( .A1(\regs[1][14] ), .A2(n998), .A3(\regs[26][14] ), .A4(
        n1002), .Y(n1407) );
  NOR4X1_LVT U1589 ( .A1(n1410), .A2(n1409), .A3(n1408), .A4(n1407), .Y(n1416)
         );
  AO22X1_LVT U1590 ( .A1(\regs[5][14] ), .A2(n987), .A3(\regs[20][14] ), .A4(
        n1001), .Y(n1414) );
  AO22X1_LVT U1591 ( .A1(\regs[13][14] ), .A2(n1025), .A3(\regs[30][14] ), 
        .A4(n975), .Y(n1413) );
  AO22X1_LVT U1592 ( .A1(\regs[29][14] ), .A2(n973), .A3(\regs[11][14] ), .A4(
        n1022), .Y(n1412) );
  AO22X1_LVT U1593 ( .A1(\regs[17][14] ), .A2(n990), .A3(\regs[16][14] ), .A4(
        n1003), .Y(n1411) );
  NOR4X1_LVT U1594 ( .A1(n1414), .A2(n1413), .A3(n1412), .A4(n1411), .Y(n1415)
         );
  NAND3X0_LVT U1595 ( .A1(n1417), .A2(n1416), .A3(n1415), .Y(n1418) );
  OR3X1_LVT U1596 ( .A1(n1420), .A2(n1419), .A3(n1418), .Y(n1421) );
  AO22X1_LVT U1597 ( .A1(wdata[14]), .A2(n960), .A3(n963), .A4(n1421), .Y(
        rdata1[14]) );
  AO22X1_LVT U1601 ( .A1(\regs[1][15] ), .A2(n998), .A3(\regs[5][15] ), .A4(
        n987), .Y(n1448) );
  AO22X1_LVT U1602 ( .A1(\regs[4][15] ), .A2(n1012), .A3(\regs[19][15] ), .A4(
        n1017), .Y(n1424) );
  INVX1_LVT U1603 ( .A(n1424), .Y(n1428) );
  AO22X1_LVT U1604 ( .A1(\regs[8][15] ), .A2(n981), .A3(\regs[16][15] ), .A4(
        n1003), .Y(n1425) );
  INVX1_LVT U1605 ( .A(n1425), .Y(n1427) );
  NAND2X0_LVT U1606 ( .A1(\regs[30][15] ), .A2(n975), .Y(n1426) );
  NAND3X0_LVT U1607 ( .A1(n1428), .A2(n1427), .A3(n1426), .Y(n1447) );
  AO22X1_LVT U1608 ( .A1(\regs[20][15] ), .A2(n1001), .A3(\regs[14][15] ), 
        .A4(n997), .Y(n1432) );
  AO22X1_LVT U1609 ( .A1(\regs[28][15] ), .A2(n986), .A3(\regs[17][15] ), .A4(
        n990), .Y(n1431) );
  AO22X1_LVT U1610 ( .A1(\regs[31][15] ), .A2(n1027), .A3(\regs[6][15] ), .A4(
        n1020), .Y(n1430) );
  AO22X1_LVT U1611 ( .A1(\regs[25][15] ), .A2(n979), .A3(\regs[3][15] ), .A4(
        n965), .Y(n1429) );
  NOR4X1_LVT U1612 ( .A1(n1432), .A2(n1431), .A3(n1430), .A4(n1429), .Y(n1445)
         );
  AO22X1_LVT U1613 ( .A1(\regs[2][15] ), .A2(n1014), .A3(\regs[27][15] ), .A4(
        n982), .Y(n1436) );
  AO22X1_LVT U1614 ( .A1(\regs[18][15] ), .A2(n995), .A3(\regs[21][15] ), .A4(
        n969), .Y(n1435) );
  AO22X1_LVT U1615 ( .A1(\regs[11][15] ), .A2(n1022), .A3(\regs[7][15] ), .A4(
        n985), .Y(n1434) );
  AO22X1_LVT U1616 ( .A1(\regs[26][15] ), .A2(n1002), .A3(\regs[9][15] ), .A4(
        n967), .Y(n1433) );
  NOR4X1_LVT U1617 ( .A1(n1436), .A2(n1435), .A3(n1434), .A4(n1433), .Y(n1444)
         );
  AO22X1_LVT U1619 ( .A1(\regs[29][15] ), .A2(n973), .A3(\regs[15][15] ), .A4(
        n1015), .Y(n1442) );
  AO22X1_LVT U1620 ( .A1(\regs[13][15] ), .A2(n1025), .A3(\regs[22][15] ), 
        .A4(n996), .Y(n1441) );
  AO22X1_LVT U1621 ( .A1(\regs[23][15] ), .A2(n968), .A3(\regs[12][15] ), .A4(
        n983), .Y(n1440) );
  AO22X1_LVT U1622 ( .A1(\regs[10][15] ), .A2(n972), .A3(\regs[24][15] ), .A4(
        n1005), .Y(n1439) );
  NOR4X1_LVT U1623 ( .A1(n1442), .A2(n1441), .A3(n1440), .A4(n1439), .Y(n1443)
         );
  NAND3X0_LVT U1624 ( .A1(n1445), .A2(n1444), .A3(n1443), .Y(n1446) );
  OR3X1_LVT U1625 ( .A1(n1448), .A2(n1447), .A3(n1446), .Y(n1449) );
  AO22X1_LVT U1626 ( .A1(wdata[15]), .A2(n960), .A3(n963), .A4(n1449), .Y(
        rdata1[15]) );
  AO22X1_LVT U1628 ( .A1(\regs[29][16] ), .A2(n973), .A3(\regs[30][16] ), .A4(
        n975), .Y(n1472) );
  AO22X1_LVT U1629 ( .A1(\regs[19][16] ), .A2(n1017), .A3(\regs[28][16] ), 
        .A4(n986), .Y(n1450) );
  INVX1_LVT U1630 ( .A(n1450), .Y(n1454) );
  AO22X1_LVT U1631 ( .A1(\regs[1][16] ), .A2(n998), .A3(\regs[12][16] ), .A4(
        n983), .Y(n1451) );
  INVX1_LVT U1632 ( .A(n1451), .Y(n1453) );
  NAND2X0_LVT U1633 ( .A1(\regs[31][16] ), .A2(n1027), .Y(n1452) );
  NAND3X0_LVT U1634 ( .A1(n1454), .A2(n1453), .A3(n1452), .Y(n1471) );
  AO22X1_LVT U1635 ( .A1(\regs[17][16] ), .A2(n990), .A3(\regs[3][16] ), .A4(
        n965), .Y(n1458) );
  AO22X1_LVT U1636 ( .A1(\regs[16][16] ), .A2(n1003), .A3(\regs[6][16] ), .A4(
        n1020), .Y(n1457) );
  AO22X1_LVT U1637 ( .A1(\regs[11][16] ), .A2(n1022), .A3(\regs[27][16] ), 
        .A4(n982), .Y(n1456) );
  AO22X1_LVT U1638 ( .A1(\regs[23][16] ), .A2(n968), .A3(\regs[15][16] ), .A4(
        n1015), .Y(n1455) );
  NOR4X1_LVT U1639 ( .A1(n1458), .A2(n1457), .A3(n1456), .A4(n1455), .Y(n1469)
         );
  AO22X1_LVT U1640 ( .A1(\regs[22][16] ), .A2(n996), .A3(\regs[21][16] ), .A4(
        n969), .Y(n1462) );
  AO22X1_LVT U1641 ( .A1(\regs[2][16] ), .A2(n1014), .A3(\regs[4][16] ), .A4(
        n1012), .Y(n1461) );
  AO22X1_LVT U1642 ( .A1(\regs[14][16] ), .A2(n997), .A3(\regs[5][16] ), .A4(
        n987), .Y(n1460) );
  AO22X1_LVT U1643 ( .A1(\regs[9][16] ), .A2(n967), .A3(\regs[20][16] ), .A4(
        n1001), .Y(n1459) );
  NOR4X1_LVT U1644 ( .A1(n1462), .A2(n1461), .A3(n1460), .A4(n1459), .Y(n1468)
         );
  AO22X1_LVT U1645 ( .A1(\regs[24][16] ), .A2(n1005), .A3(\regs[13][16] ), 
        .A4(n1025), .Y(n1466) );
  AO22X1_LVT U1646 ( .A1(\regs[26][16] ), .A2(n1002), .A3(\regs[25][16] ), 
        .A4(n979), .Y(n1465) );
  AO22X1_LVT U1647 ( .A1(\regs[18][16] ), .A2(n995), .A3(\regs[7][16] ), .A4(
        n985), .Y(n1464) );
  AO22X1_LVT U1648 ( .A1(\regs[8][16] ), .A2(n981), .A3(\regs[10][16] ), .A4(
        n972), .Y(n1463) );
  NOR4X1_LVT U1649 ( .A1(n1466), .A2(n1465), .A3(n1464), .A4(n1463), .Y(n1467)
         );
  NAND3X0_LVT U1650 ( .A1(n1469), .A2(n1468), .A3(n1467), .Y(n1470) );
  OR3X1_LVT U1651 ( .A1(n1472), .A2(n1471), .A3(n1470), .Y(n1473) );
  AO22X1_LVT U1652 ( .A1(wdata[16]), .A2(n960), .A3(n963), .A4(n1473), .Y(
        rdata1[16]) );
  AO22X1_LVT U1654 ( .A1(\regs[9][17] ), .A2(n967), .A3(\regs[27][17] ), .A4(
        n982), .Y(n1496) );
  AO22X1_LVT U1655 ( .A1(\regs[15][17] ), .A2(n1015), .A3(\regs[23][17] ), 
        .A4(n968), .Y(n1474) );
  INVX1_LVT U1656 ( .A(n1474), .Y(n1478) );
  AO22X1_LVT U1657 ( .A1(\regs[17][17] ), .A2(n990), .A3(\regs[3][17] ), .A4(
        n965), .Y(n1475) );
  INVX1_LVT U1658 ( .A(n1475), .Y(n1477) );
  NAND2X0_LVT U1659 ( .A1(\regs[20][17] ), .A2(n1001), .Y(n1476) );
  NAND3X0_LVT U1660 ( .A1(n1478), .A2(n1477), .A3(n1476), .Y(n1495) );
  AO22X1_LVT U1661 ( .A1(\regs[18][17] ), .A2(n995), .A3(\regs[14][17] ), .A4(
        n997), .Y(n1482) );
  AO22X1_LVT U1662 ( .A1(\regs[12][17] ), .A2(n983), .A3(\regs[26][17] ), .A4(
        n1002), .Y(n1481) );
  AO22X1_LVT U1663 ( .A1(\regs[6][17] ), .A2(n1020), .A3(\regs[22][17] ), .A4(
        n996), .Y(n1480) );
  AO22X1_LVT U1664 ( .A1(\regs[11][17] ), .A2(n1022), .A3(\regs[5][17] ), .A4(
        n987), .Y(n1479) );
  NOR4X1_LVT U1665 ( .A1(n1482), .A2(n1481), .A3(n1480), .A4(n1479), .Y(n1493)
         );
  AO22X1_LVT U1666 ( .A1(\regs[13][17] ), .A2(n1025), .A3(\regs[10][17] ), 
        .A4(n972), .Y(n1486) );
  AO22X1_LVT U1667 ( .A1(\regs[31][17] ), .A2(n1027), .A3(\regs[8][17] ), .A4(
        n981), .Y(n1485) );
  AO22X1_LVT U1668 ( .A1(\regs[1][17] ), .A2(n998), .A3(\regs[19][17] ), .A4(
        n1017), .Y(n1484) );
  AO22X1_LVT U1669 ( .A1(\regs[30][17] ), .A2(n975), .A3(\regs[29][17] ), .A4(
        n973), .Y(n1483) );
  NOR4X1_LVT U1670 ( .A1(n1486), .A2(n1485), .A3(n1484), .A4(n1483), .Y(n1492)
         );
  AO22X1_LVT U1671 ( .A1(\regs[4][17] ), .A2(n1012), .A3(\regs[7][17] ), .A4(
        n985), .Y(n1490) );
  AO22X1_LVT U1672 ( .A1(\regs[2][17] ), .A2(n1014), .A3(\regs[28][17] ), .A4(
        n986), .Y(n1489) );
  AO22X1_LVT U1673 ( .A1(\regs[16][17] ), .A2(n1003), .A3(\regs[25][17] ), 
        .A4(n979), .Y(n1488) );
  AO22X1_LVT U1674 ( .A1(\regs[24][17] ), .A2(n1005), .A3(\regs[21][17] ), 
        .A4(n969), .Y(n1487) );
  NOR4X1_LVT U1675 ( .A1(n1490), .A2(n1489), .A3(n1488), .A4(n1487), .Y(n1491)
         );
  NAND3X0_LVT U1676 ( .A1(n1493), .A2(n1492), .A3(n1491), .Y(n1494) );
  OR3X1_LVT U1677 ( .A1(n1496), .A2(n1495), .A3(n1494), .Y(n1497) );
  AO22X1_LVT U1678 ( .A1(wdata[17]), .A2(n960), .A3(n963), .A4(n1497), .Y(
        rdata1[17]) );
  AO22X1_LVT U1680 ( .A1(\regs[11][18] ), .A2(n1022), .A3(\regs[8][18] ), .A4(
        n981), .Y(n1520) );
  AO22X1_LVT U1681 ( .A1(\regs[20][18] ), .A2(n1001), .A3(\regs[9][18] ), .A4(
        n967), .Y(n1498) );
  INVX1_LVT U1682 ( .A(n1498), .Y(n1502) );
  AO22X1_LVT U1683 ( .A1(\regs[25][18] ), .A2(n979), .A3(\regs[18][18] ), .A4(
        n995), .Y(n1499) );
  INVX1_LVT U1684 ( .A(n1499), .Y(n1501) );
  NAND2X0_LVT U1685 ( .A1(\regs[7][18] ), .A2(n985), .Y(n1500) );
  NAND3X0_LVT U1686 ( .A1(n1502), .A2(n1501), .A3(n1500), .Y(n1519) );
  AO22X1_LVT U1687 ( .A1(\regs[30][18] ), .A2(n975), .A3(\regs[24][18] ), .A4(
        n1005), .Y(n1506) );
  AO22X1_LVT U1688 ( .A1(\regs[31][18] ), .A2(n1027), .A3(\regs[13][18] ), 
        .A4(n1025), .Y(n1505) );
  AO22X1_LVT U1689 ( .A1(\regs[21][18] ), .A2(n969), .A3(\regs[26][18] ), .A4(
        n1002), .Y(n1504) );
  AO22X1_LVT U1690 ( .A1(\regs[22][18] ), .A2(n996), .A3(\regs[1][18] ), .A4(
        n998), .Y(n1503) );
  NOR4X1_LVT U1691 ( .A1(n1506), .A2(n1505), .A3(n1504), .A4(n1503), .Y(n1517)
         );
  AO22X1_LVT U1692 ( .A1(\regs[27][18] ), .A2(n982), .A3(\regs[5][18] ), .A4(
        n987), .Y(n1510) );
  AO22X1_LVT U1693 ( .A1(\regs[17][18] ), .A2(n990), .A3(\regs[15][18] ), .A4(
        n1015), .Y(n1509) );
  AO22X1_LVT U1694 ( .A1(\regs[4][18] ), .A2(n1012), .A3(\regs[6][18] ), .A4(
        n1020), .Y(n1508) );
  AO22X1_LVT U1695 ( .A1(\regs[23][18] ), .A2(n968), .A3(\regs[10][18] ), .A4(
        n972), .Y(n1507) );
  NOR4X1_LVT U1696 ( .A1(n1510), .A2(n1509), .A3(n1508), .A4(n1507), .Y(n1516)
         );
  AO22X1_LVT U1697 ( .A1(\regs[14][18] ), .A2(n997), .A3(\regs[28][18] ), .A4(
        n986), .Y(n1514) );
  AO22X1_LVT U1698 ( .A1(\regs[2][18] ), .A2(n1014), .A3(\regs[12][18] ), .A4(
        n983), .Y(n1513) );
  AO22X1_LVT U1699 ( .A1(\regs[16][18] ), .A2(n1003), .A3(\regs[29][18] ), 
        .A4(n973), .Y(n1512) );
  AO22X1_LVT U1700 ( .A1(\regs[3][18] ), .A2(n965), .A3(\regs[19][18] ), .A4(
        n1017), .Y(n1511) );
  NOR4X1_LVT U1701 ( .A1(n1514), .A2(n1513), .A3(n1512), .A4(n1511), .Y(n1515)
         );
  NAND3X0_LVT U1702 ( .A1(n1517), .A2(n1516), .A3(n1515), .Y(n1518) );
  OR3X1_LVT U1703 ( .A1(n1520), .A2(n1519), .A3(n1518), .Y(n1521) );
  AO22X1_LVT U1704 ( .A1(wdata[18]), .A2(n960), .A3(n963), .A4(n1521), .Y(
        rdata1[18]) );
  AO22X1_LVT U1706 ( .A1(\regs[2][19] ), .A2(n1014), .A3(\regs[12][19] ), .A4(
        n983), .Y(n2536) );
  AO22X1_LVT U1707 ( .A1(\regs[22][19] ), .A2(n996), .A3(\regs[26][19] ), .A4(
        n1002), .Y(n1522) );
  INVX1_LVT U1708 ( .A(n1522), .Y(n1526) );
  AO22X1_LVT U1709 ( .A1(\regs[7][19] ), .A2(n985), .A3(\regs[17][19] ), .A4(
        n990), .Y(n1523) );
  INVX1_LVT U1710 ( .A(n1523), .Y(n1525) );
  NAND2X0_LVT U1711 ( .A1(\regs[28][19] ), .A2(n986), .Y(n1524) );
  NAND3X0_LVT U1712 ( .A1(n1526), .A2(n1525), .A3(n1524), .Y(n2535) );
  AO22X1_LVT U1713 ( .A1(\regs[18][19] ), .A2(n995), .A3(\regs[14][19] ), .A4(
        n997), .Y(n1530) );
  AO22X1_LVT U1714 ( .A1(\regs[19][19] ), .A2(n1017), .A3(\regs[31][19] ), 
        .A4(n1027), .Y(n1529) );
  AO22X1_LVT U1715 ( .A1(\regs[23][19] ), .A2(n968), .A3(\regs[3][19] ), .A4(
        n965), .Y(n1528) );
  AO22X1_LVT U1716 ( .A1(\regs[9][19] ), .A2(n967), .A3(\regs[6][19] ), .A4(
        n1020), .Y(n1527) );
  NOR4X1_LVT U1717 ( .A1(n1530), .A2(n1529), .A3(n1528), .A4(n1527), .Y(n2533)
         );
  AO22X1_LVT U1718 ( .A1(\regs[24][19] ), .A2(n1005), .A3(\regs[25][19] ), 
        .A4(n979), .Y(n1534) );
  AO22X1_LVT U1719 ( .A1(\regs[30][19] ), .A2(n975), .A3(\regs[10][19] ), .A4(
        n972), .Y(n1533) );
  AO22X1_LVT U1720 ( .A1(\regs[1][19] ), .A2(n998), .A3(\regs[15][19] ), .A4(
        n1015), .Y(n1532) );
  AO22X1_LVT U1721 ( .A1(\regs[20][19] ), .A2(n1001), .A3(\regs[16][19] ), 
        .A4(n1003), .Y(n1531) );
  NOR4X1_LVT U1722 ( .A1(n1534), .A2(n1533), .A3(n1532), .A4(n1531), .Y(n2532)
         );
  AO22X1_LVT U1723 ( .A1(\regs[29][19] ), .A2(n973), .A3(\regs[8][19] ), .A4(
        n981), .Y(n1538) );
  AO22X1_LVT U1724 ( .A1(\regs[11][19] ), .A2(n1022), .A3(\regs[5][19] ), .A4(
        n987), .Y(n1537) );
  AO22X1_LVT U1725 ( .A1(\regs[27][19] ), .A2(n982), .A3(\regs[13][19] ), .A4(
        n1025), .Y(n1536) );
  AO22X1_LVT U1726 ( .A1(\regs[4][19] ), .A2(n1012), .A3(\regs[21][19] ), .A4(
        n969), .Y(n1535) );
  NOR4X1_LVT U1727 ( .A1(n1538), .A2(n1537), .A3(n1536), .A4(n1535), .Y(n2531)
         );
  NAND3X0_LVT U1728 ( .A1(n2533), .A2(n2532), .A3(n2531), .Y(n2534) );
  OR3X1_LVT U1729 ( .A1(n2536), .A2(n2535), .A3(n2534), .Y(n2537) );
  AO22X1_LVT U1730 ( .A1(wdata[19]), .A2(n960), .A3(n963), .A4(n2537), .Y(
        rdata1[19]) );
  AO22X1_LVT U1732 ( .A1(\regs[9][20] ), .A2(n967), .A3(\regs[18][20] ), .A4(
        n995), .Y(n2560) );
  AO22X1_LVT U1733 ( .A1(\regs[4][20] ), .A2(n1012), .A3(\regs[11][20] ), .A4(
        n1022), .Y(n2538) );
  INVX1_LVT U1734 ( .A(n2538), .Y(n2542) );
  AO22X1_LVT U1735 ( .A1(\regs[2][20] ), .A2(n1014), .A3(\regs[3][20] ), .A4(
        n965), .Y(n2539) );
  INVX1_LVT U1736 ( .A(n2539), .Y(n2541) );
  NAND2X0_LVT U1737 ( .A1(\regs[16][20] ), .A2(n1003), .Y(n2540) );
  NAND3X0_LVT U1738 ( .A1(n2542), .A2(n2541), .A3(n2540), .Y(n2559) );
  AO22X1_LVT U1739 ( .A1(\regs[10][20] ), .A2(n972), .A3(\regs[17][20] ), .A4(
        n990), .Y(n2546) );
  AO22X1_LVT U1740 ( .A1(\regs[13][20] ), .A2(n1025), .A3(\regs[6][20] ), .A4(
        n1020), .Y(n2545) );
  AO22X1_LVT U1741 ( .A1(\regs[14][20] ), .A2(n997), .A3(\regs[24][20] ), .A4(
        n1005), .Y(n2544) );
  AO22X1_LVT U1742 ( .A1(\regs[7][20] ), .A2(n985), .A3(\regs[8][20] ), .A4(
        n981), .Y(n2543) );
  NOR4X1_LVT U1743 ( .A1(n2546), .A2(n2545), .A3(n2544), .A4(n2543), .Y(n2557)
         );
  AO22X1_LVT U1744 ( .A1(\regs[20][20] ), .A2(n1001), .A3(\regs[12][20] ), 
        .A4(n983), .Y(n2550) );
  AO22X1_LVT U1745 ( .A1(\regs[27][20] ), .A2(n982), .A3(\regs[21][20] ), .A4(
        n969), .Y(n2549) );
  AO22X1_LVT U1746 ( .A1(\regs[25][20] ), .A2(n979), .A3(\regs[29][20] ), .A4(
        n973), .Y(n2548) );
  AO22X1_LVT U1747 ( .A1(\regs[28][20] ), .A2(n986), .A3(\regs[22][20] ), .A4(
        n996), .Y(n2547) );
  NOR4X1_LVT U1748 ( .A1(n2550), .A2(n2549), .A3(n2548), .A4(n2547), .Y(n2556)
         );
  AO22X1_LVT U1749 ( .A1(\regs[1][20] ), .A2(n998), .A3(\regs[5][20] ), .A4(
        n987), .Y(n2554) );
  AO22X1_LVT U1750 ( .A1(\regs[19][20] ), .A2(n1017), .A3(\regs[31][20] ), 
        .A4(n1027), .Y(n2553) );
  AO22X1_LVT U1751 ( .A1(\regs[15][20] ), .A2(n1015), .A3(\regs[23][20] ), 
        .A4(n968), .Y(n2552) );
  AO22X1_LVT U1752 ( .A1(\regs[26][20] ), .A2(n1002), .A3(\regs[30][20] ), 
        .A4(n975), .Y(n2551) );
  NOR4X1_LVT U1753 ( .A1(n2554), .A2(n2553), .A3(n2552), .A4(n2551), .Y(n2555)
         );
  NAND3X0_LVT U1754 ( .A1(n2557), .A2(n2556), .A3(n2555), .Y(n2558) );
  OR3X1_LVT U1755 ( .A1(n2560), .A2(n2559), .A3(n2558), .Y(n2561) );
  AO22X1_LVT U1756 ( .A1(wdata[20]), .A2(n960), .A3(n963), .A4(n2561), .Y(
        rdata1[20]) );
  AO22X1_LVT U1758 ( .A1(\regs[4][21] ), .A2(n1012), .A3(\regs[9][21] ), .A4(
        n967), .Y(n2584) );
  AO22X1_LVT U1759 ( .A1(\regs[29][21] ), .A2(n973), .A3(\regs[8][21] ), .A4(
        n981), .Y(n2562) );
  INVX1_LVT U1760 ( .A(n2562), .Y(n2566) );
  AO22X1_LVT U1761 ( .A1(\regs[7][21] ), .A2(n985), .A3(\regs[26][21] ), .A4(
        n1002), .Y(n2563) );
  INVX1_LVT U1762 ( .A(n2563), .Y(n2565) );
  NAND2X0_LVT U1763 ( .A1(\regs[19][21] ), .A2(n1017), .Y(n2564) );
  NAND3X0_LVT U1764 ( .A1(n2566), .A2(n2565), .A3(n2564), .Y(n2583) );
  AO22X1_LVT U1765 ( .A1(\regs[14][21] ), .A2(n997), .A3(\regs[10][21] ), .A4(
        n972), .Y(n2570) );
  AO22X1_LVT U1766 ( .A1(\regs[27][21] ), .A2(n982), .A3(\regs[18][21] ), .A4(
        n995), .Y(n2569) );
  AO22X1_LVT U1767 ( .A1(\regs[12][21] ), .A2(n983), .A3(\regs[31][21] ), .A4(
        n1027), .Y(n2568) );
  AO22X1_LVT U1768 ( .A1(\regs[23][21] ), .A2(n968), .A3(\regs[1][21] ), .A4(
        n998), .Y(n2567) );
  NOR4X1_LVT U1769 ( .A1(n2570), .A2(n2569), .A3(n2568), .A4(n2567), .Y(n2581)
         );
  AO22X1_LVT U1770 ( .A1(\regs[6][21] ), .A2(n1020), .A3(\regs[22][21] ), .A4(
        n996), .Y(n2574) );
  AO22X1_LVT U1771 ( .A1(\regs[20][21] ), .A2(n1001), .A3(\regs[25][21] ), 
        .A4(n979), .Y(n2573) );
  AO22X1_LVT U1772 ( .A1(\regs[13][21] ), .A2(n1025), .A3(\regs[21][21] ), 
        .A4(n969), .Y(n2572) );
  AO22X1_LVT U1773 ( .A1(\regs[16][21] ), .A2(n1003), .A3(\regs[3][21] ), .A4(
        n965), .Y(n2571) );
  NOR4X1_LVT U1774 ( .A1(n2574), .A2(n2573), .A3(n2572), .A4(n2571), .Y(n2580)
         );
  AO22X1_LVT U1775 ( .A1(\regs[11][21] ), .A2(n1022), .A3(\regs[17][21] ), 
        .A4(n990), .Y(n2578) );
  AO22X1_LVT U1776 ( .A1(\regs[15][21] ), .A2(n1015), .A3(\regs[28][21] ), 
        .A4(n986), .Y(n2577) );
  AO22X1_LVT U1777 ( .A1(\regs[24][21] ), .A2(n1005), .A3(\regs[5][21] ), .A4(
        n987), .Y(n2576) );
  AO22X1_LVT U1778 ( .A1(\regs[30][21] ), .A2(n975), .A3(\regs[2][21] ), .A4(
        n1014), .Y(n2575) );
  NOR4X1_LVT U1779 ( .A1(n2578), .A2(n2577), .A3(n2576), .A4(n2575), .Y(n2579)
         );
  NAND3X0_LVT U1780 ( .A1(n2581), .A2(n2580), .A3(n2579), .Y(n2582) );
  OR3X1_LVT U1781 ( .A1(n2584), .A2(n2583), .A3(n2582), .Y(n2585) );
  AO22X1_LVT U1782 ( .A1(wdata[21]), .A2(n960), .A3(n963), .A4(n2585), .Y(
        rdata1[21]) );
  AO22X1_LVT U1784 ( .A1(\regs[29][22] ), .A2(n973), .A3(\regs[20][22] ), .A4(
        n1001), .Y(n2610) );
  AO22X1_LVT U1786 ( .A1(\regs[31][22] ), .A2(n1027), .A3(\regs[27][22] ), 
        .A4(n982), .Y(n2588) );
  INVX1_LVT U1787 ( .A(n2588), .Y(n2592) );
  AO22X1_LVT U1788 ( .A1(\regs[21][22] ), .A2(n969), .A3(\regs[15][22] ), .A4(
        n1015), .Y(n2589) );
  INVX1_LVT U1789 ( .A(n2589), .Y(n2591) );
  NAND2X0_LVT U1790 ( .A1(\regs[30][22] ), .A2(n975), .Y(n2590) );
  NAND3X0_LVT U1791 ( .A1(n2592), .A2(n2591), .A3(n2590), .Y(n2609) );
  AO22X1_LVT U1792 ( .A1(\regs[18][22] ), .A2(n995), .A3(\regs[19][22] ), .A4(
        n1017), .Y(n2596) );
  AO22X1_LVT U1793 ( .A1(\regs[3][22] ), .A2(n965), .A3(\regs[24][22] ), .A4(
        n1005), .Y(n2595) );
  AO22X1_LVT U1794 ( .A1(\regs[17][22] ), .A2(n990), .A3(\regs[28][22] ), .A4(
        n986), .Y(n2594) );
  AO22X1_LVT U1795 ( .A1(\regs[9][22] ), .A2(n967), .A3(\regs[13][22] ), .A4(
        n1025), .Y(n2593) );
  NOR4X1_LVT U1796 ( .A1(n2596), .A2(n2595), .A3(n2594), .A4(n2593), .Y(n2607)
         );
  AO22X1_LVT U1797 ( .A1(\regs[14][22] ), .A2(n997), .A3(\regs[12][22] ), .A4(
        n983), .Y(n2600) );
  AO22X1_LVT U1798 ( .A1(\regs[2][22] ), .A2(n1014), .A3(\regs[4][22] ), .A4(
        n1012), .Y(n2599) );
  AO22X1_LVT U1799 ( .A1(\regs[16][22] ), .A2(n1003), .A3(\regs[7][22] ), .A4(
        n985), .Y(n2598) );
  AO22X1_LVT U1800 ( .A1(\regs[5][22] ), .A2(n987), .A3(\regs[6][22] ), .A4(
        n1020), .Y(n2597) );
  NOR4X1_LVT U1801 ( .A1(n2600), .A2(n2599), .A3(n2598), .A4(n2597), .Y(n2606)
         );
  AO22X1_LVT U1802 ( .A1(\regs[25][22] ), .A2(n979), .A3(\regs[8][22] ), .A4(
        n981), .Y(n2604) );
  AO22X1_LVT U1803 ( .A1(\regs[1][22] ), .A2(n998), .A3(\regs[22][22] ), .A4(
        n996), .Y(n2603) );
  AO22X1_LVT U1804 ( .A1(\regs[10][22] ), .A2(n972), .A3(\regs[23][22] ), .A4(
        n968), .Y(n2602) );
  AO22X1_LVT U1805 ( .A1(\regs[11][22] ), .A2(n1022), .A3(\regs[26][22] ), 
        .A4(n1002), .Y(n2601) );
  NOR4X1_LVT U1806 ( .A1(n2604), .A2(n2603), .A3(n2602), .A4(n2601), .Y(n2605)
         );
  NAND3X0_LVT U1807 ( .A1(n2607), .A2(n2606), .A3(n2605), .Y(n2608) );
  OR3X1_LVT U1808 ( .A1(n2610), .A2(n2609), .A3(n2608), .Y(n2611) );
  AO22X1_LVT U1809 ( .A1(wdata[22]), .A2(n960), .A3(n963), .A4(n2611), .Y(
        rdata1[22]) );
  AO22X1_LVT U1811 ( .A1(\regs[4][23] ), .A2(n1012), .A3(\regs[23][23] ), .A4(
        n968), .Y(n2634) );
  AO22X1_LVT U1812 ( .A1(\regs[6][23] ), .A2(n1020), .A3(\regs[25][23] ), .A4(
        n979), .Y(n2612) );
  INVX1_LVT U1813 ( .A(n2612), .Y(n2616) );
  AO22X1_LVT U1814 ( .A1(\regs[10][23] ), .A2(n972), .A3(\regs[20][23] ), .A4(
        n1001), .Y(n2613) );
  INVX1_LVT U1815 ( .A(n2613), .Y(n2615) );
  NAND2X0_LVT U1816 ( .A1(\regs[7][23] ), .A2(n985), .Y(n2614) );
  NAND3X0_LVT U1817 ( .A1(n2616), .A2(n2615), .A3(n2614), .Y(n2633) );
  AO22X1_LVT U1818 ( .A1(\regs[5][23] ), .A2(n987), .A3(\regs[12][23] ), .A4(
        n983), .Y(n2620) );
  AO22X1_LVT U1819 ( .A1(\regs[18][23] ), .A2(n995), .A3(\regs[24][23] ), .A4(
        n1005), .Y(n2619) );
  AO22X1_LVT U1820 ( .A1(\regs[1][23] ), .A2(n998), .A3(\regs[17][23] ), .A4(
        n990), .Y(n2618) );
  AO22X1_LVT U1821 ( .A1(\regs[16][23] ), .A2(n1003), .A3(\regs[26][23] ), 
        .A4(n1002), .Y(n2617) );
  NOR4X1_LVT U1822 ( .A1(n2620), .A2(n2619), .A3(n2618), .A4(n2617), .Y(n2631)
         );
  AO22X1_LVT U1823 ( .A1(\regs[19][23] ), .A2(n1017), .A3(\regs[28][23] ), 
        .A4(n986), .Y(n2624) );
  AO22X1_LVT U1824 ( .A1(\regs[13][23] ), .A2(n1025), .A3(\regs[8][23] ), .A4(
        n981), .Y(n2623) );
  AO22X1_LVT U1825 ( .A1(\regs[9][23] ), .A2(n967), .A3(\regs[3][23] ), .A4(
        n965), .Y(n2622) );
  AO22X1_LVT U1826 ( .A1(\regs[15][23] ), .A2(n1015), .A3(\regs[27][23] ), 
        .A4(n982), .Y(n2621) );
  NOR4X1_LVT U1827 ( .A1(n2624), .A2(n2623), .A3(n2622), .A4(n2621), .Y(n2630)
         );
  AO22X1_LVT U1828 ( .A1(\regs[22][23] ), .A2(n996), .A3(\regs[29][23] ), .A4(
        n973), .Y(n2628) );
  AO22X1_LVT U1829 ( .A1(\regs[2][23] ), .A2(n1014), .A3(\regs[31][23] ), .A4(
        n1027), .Y(n2627) );
  AO22X1_LVT U1830 ( .A1(\regs[21][23] ), .A2(n969), .A3(\regs[30][23] ), .A4(
        n975), .Y(n2626) );
  AO22X1_LVT U1831 ( .A1(\regs[11][23] ), .A2(n1022), .A3(\regs[14][23] ), 
        .A4(n997), .Y(n2625) );
  NOR4X1_LVT U1832 ( .A1(n2628), .A2(n2627), .A3(n2626), .A4(n2625), .Y(n2629)
         );
  NAND3X0_LVT U1833 ( .A1(n2631), .A2(n2630), .A3(n2629), .Y(n2632) );
  OR3X1_LVT U1834 ( .A1(n2634), .A2(n2633), .A3(n2632), .Y(n2635) );
  AO22X1_LVT U1835 ( .A1(wdata[23]), .A2(n960), .A3(n963), .A4(n2635), .Y(
        rdata1[23]) );
  AO22X1_LVT U1837 ( .A1(\regs[2][24] ), .A2(n1014), .A3(\regs[14][24] ), .A4(
        n997), .Y(n2659) );
  AO22X1_LVT U1838 ( .A1(\regs[20][24] ), .A2(n1001), .A3(\regs[4][24] ), .A4(
        n1012), .Y(n2637) );
  INVX1_LVT U1839 ( .A(n2637), .Y(n2641) );
  AO22X1_LVT U1840 ( .A1(\regs[25][24] ), .A2(n979), .A3(\regs[23][24] ), .A4(
        n968), .Y(n2638) );
  INVX1_LVT U1841 ( .A(n2638), .Y(n2640) );
  NAND2X0_LVT U1842 ( .A1(\regs[13][24] ), .A2(n1025), .Y(n2639) );
  NAND3X0_LVT U1843 ( .A1(n2641), .A2(n2640), .A3(n2639), .Y(n2658) );
  AO22X1_LVT U1844 ( .A1(\regs[1][24] ), .A2(n998), .A3(\regs[30][24] ), .A4(
        n975), .Y(n2645) );
  AO22X1_LVT U1845 ( .A1(\regs[27][24] ), .A2(n982), .A3(\regs[22][24] ), .A4(
        n996), .Y(n2644) );
  AO22X1_LVT U1846 ( .A1(\regs[24][24] ), .A2(n1005), .A3(\regs[26][24] ), 
        .A4(n1002), .Y(n2643) );
  AO22X1_LVT U1847 ( .A1(\regs[5][24] ), .A2(n987), .A3(\regs[28][24] ), .A4(
        n986), .Y(n2642) );
  NOR4X1_LVT U1848 ( .A1(n2645), .A2(n2644), .A3(n2643), .A4(n2642), .Y(n2656)
         );
  AO22X1_LVT U1849 ( .A1(\regs[9][24] ), .A2(n967), .A3(\regs[8][24] ), .A4(
        n981), .Y(n2649) );
  AO22X1_LVT U1850 ( .A1(\regs[11][24] ), .A2(n1022), .A3(\regs[29][24] ), 
        .A4(n973), .Y(n2648) );
  AO22X1_LVT U1851 ( .A1(\regs[21][24] ), .A2(n969), .A3(\regs[15][24] ), .A4(
        n1015), .Y(n2647) );
  AO22X1_LVT U1852 ( .A1(\regs[18][24] ), .A2(n995), .A3(\regs[3][24] ), .A4(
        n965), .Y(n2646) );
  NOR4X1_LVT U1853 ( .A1(n2649), .A2(n2648), .A3(n2647), .A4(n2646), .Y(n2655)
         );
  AO22X1_LVT U1854 ( .A1(\regs[10][24] ), .A2(n972), .A3(\regs[6][24] ), .A4(
        n1020), .Y(n2653) );
  AO22X1_LVT U1855 ( .A1(\regs[16][24] ), .A2(n1003), .A3(\regs[7][24] ), .A4(
        n985), .Y(n2652) );
  AO22X1_LVT U1856 ( .A1(\regs[12][24] ), .A2(n983), .A3(\regs[31][24] ), .A4(
        n3481), .Y(n2651) );
  AO22X1_LVT U1857 ( .A1(\regs[19][24] ), .A2(n1017), .A3(\regs[17][24] ), 
        .A4(n990), .Y(n2650) );
  NOR4X1_LVT U1858 ( .A1(n2653), .A2(n2652), .A3(n2651), .A4(n2650), .Y(n2654)
         );
  NAND3X0_LVT U1859 ( .A1(n2656), .A2(n2655), .A3(n2654), .Y(n2657) );
  OR3X1_LVT U1860 ( .A1(n2659), .A2(n2658), .A3(n2657), .Y(n2660) );
  AO22X1_LVT U1861 ( .A1(wdata[24]), .A2(n960), .A3(n963), .A4(n2660), .Y(
        rdata1[24]) );
  AO22X1_LVT U1863 ( .A1(\regs[13][25] ), .A2(n1025), .A3(\regs[10][25] ), 
        .A4(n972), .Y(n2683) );
  AO22X1_LVT U1864 ( .A1(\regs[16][25] ), .A2(n1003), .A3(\regs[17][25] ), 
        .A4(n990), .Y(n2661) );
  INVX1_LVT U1865 ( .A(n2661), .Y(n2665) );
  AO22X1_LVT U1866 ( .A1(\regs[7][25] ), .A2(n985), .A3(\regs[1][25] ), .A4(
        n998), .Y(n2662) );
  INVX1_LVT U1867 ( .A(n2662), .Y(n2664) );
  NAND2X0_LVT U1868 ( .A1(\regs[5][25] ), .A2(n987), .Y(n2663) );
  NAND3X0_LVT U1869 ( .A1(n2665), .A2(n2664), .A3(n2663), .Y(n2682) );
  AO22X1_LVT U1870 ( .A1(\regs[27][25] ), .A2(n982), .A3(\regs[26][25] ), .A4(
        n1002), .Y(n2669) );
  AO22X1_LVT U1871 ( .A1(\regs[24][25] ), .A2(n1005), .A3(\regs[11][25] ), 
        .A4(n1022), .Y(n2668) );
  AO22X1_LVT U1872 ( .A1(\regs[12][25] ), .A2(n983), .A3(\regs[30][25] ), .A4(
        n975), .Y(n2667) );
  AO22X1_LVT U1873 ( .A1(\regs[14][25] ), .A2(n997), .A3(\regs[6][25] ), .A4(
        n1020), .Y(n2666) );
  NOR4X1_LVT U1874 ( .A1(n2669), .A2(n2668), .A3(n2667), .A4(n2666), .Y(n2680)
         );
  AO22X1_LVT U1875 ( .A1(\regs[25][25] ), .A2(n979), .A3(\regs[18][25] ), .A4(
        n995), .Y(n2673) );
  AO22X1_LVT U1876 ( .A1(\regs[22][25] ), .A2(n996), .A3(\regs[4][25] ), .A4(
        n1012), .Y(n2672) );
  AO22X1_LVT U1877 ( .A1(\regs[21][25] ), .A2(n3475), .A3(\regs[19][25] ), 
        .A4(n1017), .Y(n2671) );
  AO22X1_LVT U1878 ( .A1(\regs[23][25] ), .A2(n968), .A3(\regs[20][25] ), .A4(
        n1001), .Y(n2670) );
  NOR4X1_LVT U1879 ( .A1(n2673), .A2(n2672), .A3(n2671), .A4(n2670), .Y(n2679)
         );
  AO22X1_LVT U1880 ( .A1(\regs[28][25] ), .A2(n986), .A3(\regs[29][25] ), .A4(
        n973), .Y(n2677) );
  AO22X1_LVT U1881 ( .A1(\regs[9][25] ), .A2(n967), .A3(\regs[15][25] ), .A4(
        n1015), .Y(n2676) );
  AO22X1_LVT U1882 ( .A1(\regs[31][25] ), .A2(n1027), .A3(\regs[8][25] ), .A4(
        n981), .Y(n2675) );
  AO22X1_LVT U1883 ( .A1(\regs[3][25] ), .A2(n965), .A3(\regs[2][25] ), .A4(
        n1014), .Y(n2674) );
  NOR4X1_LVT U1884 ( .A1(n2677), .A2(n2676), .A3(n2675), .A4(n2674), .Y(n2678)
         );
  NAND3X0_LVT U1885 ( .A1(n2680), .A2(n2679), .A3(n2678), .Y(n2681) );
  OR3X1_LVT U1886 ( .A1(n2683), .A2(n2682), .A3(n2681), .Y(n2684) );
  AO22X1_LVT U1887 ( .A1(wdata[25]), .A2(n960), .A3(n963), .A4(n2684), .Y(
        rdata1[25]) );
  AO22X1_LVT U1889 ( .A1(\regs[12][26] ), .A2(n983), .A3(\regs[20][26] ), .A4(
        n1001), .Y(n2710) );
  AO22X1_LVT U1890 ( .A1(\regs[19][26] ), .A2(n1017), .A3(\regs[21][26] ), 
        .A4(n3475), .Y(n2685) );
  INVX1_LVT U1891 ( .A(n2685), .Y(n2691) );
  AO22X1_LVT U1892 ( .A1(\regs[30][26] ), .A2(n975), .A3(\regs[18][26] ), .A4(
        n995), .Y(n2688) );
  INVX1_LVT U1893 ( .A(n2688), .Y(n2690) );
  NAND2X0_LVT U1894 ( .A1(\regs[24][26] ), .A2(n1005), .Y(n2689) );
  NAND3X0_LVT U1895 ( .A1(n2691), .A2(n2690), .A3(n2689), .Y(n2709) );
  AO22X1_LVT U1896 ( .A1(\regs[2][26] ), .A2(n1014), .A3(\regs[6][26] ), .A4(
        n1020), .Y(n2696) );
  AO22X1_LVT U1897 ( .A1(\regs[31][26] ), .A2(n3481), .A3(\regs[3][26] ), .A4(
        n965), .Y(n2695) );
  AO22X1_LVT U1898 ( .A1(\regs[8][26] ), .A2(n981), .A3(\regs[16][26] ), .A4(
        n1003), .Y(n2694) );
  AO22X1_LVT U1899 ( .A1(\regs[28][26] ), .A2(n986), .A3(\regs[13][26] ), .A4(
        n1025), .Y(n2693) );
  NOR4X1_LVT U1900 ( .A1(n2696), .A2(n2695), .A3(n2694), .A4(n2693), .Y(n2707)
         );
  AO22X1_LVT U1901 ( .A1(\regs[15][26] ), .A2(n1015), .A3(\regs[17][26] ), 
        .A4(n990), .Y(n2700) );
  AO22X1_LVT U1902 ( .A1(\regs[23][26] ), .A2(n968), .A3(\regs[25][26] ), .A4(
        n979), .Y(n2699) );
  AO22X1_LVT U1903 ( .A1(\regs[22][26] ), .A2(n996), .A3(\regs[4][26] ), .A4(
        n1012), .Y(n2698) );
  AO22X1_LVT U1904 ( .A1(\regs[5][26] ), .A2(n987), .A3(\regs[7][26] ), .A4(
        n985), .Y(n2697) );
  NOR4X1_LVT U1905 ( .A1(n2700), .A2(n2699), .A3(n2698), .A4(n2697), .Y(n2706)
         );
  AO22X1_LVT U1906 ( .A1(\regs[11][26] ), .A2(n1022), .A3(\regs[29][26] ), 
        .A4(n973), .Y(n2704) );
  AO22X1_LVT U1907 ( .A1(\regs[14][26] ), .A2(n997), .A3(\regs[1][26] ), .A4(
        n998), .Y(n2703) );
  AO22X1_LVT U1908 ( .A1(\regs[9][26] ), .A2(n967), .A3(\regs[27][26] ), .A4(
        n982), .Y(n2702) );
  AO22X1_LVT U1909 ( .A1(\regs[10][26] ), .A2(n972), .A3(\regs[26][26] ), .A4(
        n1002), .Y(n2701) );
  NOR4X1_LVT U1910 ( .A1(n2704), .A2(n2703), .A3(n2702), .A4(n2701), .Y(n2705)
         );
  NAND3X0_LVT U1911 ( .A1(n2707), .A2(n2706), .A3(n2705), .Y(n2708) );
  OR3X1_LVT U1912 ( .A1(n2710), .A2(n2709), .A3(n2708), .Y(n2711) );
  AO22X1_LVT U1913 ( .A1(wdata[26]), .A2(n960), .A3(n963), .A4(n2711), .Y(
        rdata1[26]) );
  AO22X1_LVT U1915 ( .A1(\regs[20][27] ), .A2(n1001), .A3(\regs[28][27] ), 
        .A4(n986), .Y(n2737) );
  AO22X1_LVT U1916 ( .A1(\regs[13][27] ), .A2(n1025), .A3(\regs[11][27] ), 
        .A4(n1022), .Y(n2712) );
  INVX1_LVT U1917 ( .A(n2712), .Y(n2716) );
  AO22X1_LVT U1918 ( .A1(\regs[5][27] ), .A2(n987), .A3(\regs[25][27] ), .A4(
        n979), .Y(n2713) );
  INVX1_LVT U1919 ( .A(n2713), .Y(n2715) );
  NAND2X0_LVT U1920 ( .A1(\regs[10][27] ), .A2(n972), .Y(n2714) );
  NAND3X0_LVT U1921 ( .A1(n2716), .A2(n2715), .A3(n2714), .Y(n2736) );
  AO22X1_LVT U1922 ( .A1(\regs[23][27] ), .A2(n968), .A3(\regs[21][27] ), .A4(
        n3475), .Y(n2722) );
  AO22X1_LVT U1923 ( .A1(\regs[16][27] ), .A2(n1003), .A3(\regs[24][27] ), 
        .A4(n1005), .Y(n2721) );
  AO22X1_LVT U1924 ( .A1(\regs[15][27] ), .A2(n1015), .A3(\regs[1][27] ), .A4(
        n998), .Y(n2720) );
  AO22X1_LVT U1925 ( .A1(\regs[27][27] ), .A2(n982), .A3(\regs[4][27] ), .A4(
        n1012), .Y(n2719) );
  NOR4X1_LVT U1926 ( .A1(n2722), .A2(n2721), .A3(n2720), .A4(n2719), .Y(n2734)
         );
  AO22X1_LVT U1927 ( .A1(\regs[6][27] ), .A2(n1020), .A3(\regs[14][27] ), .A4(
        n997), .Y(n2726) );
  AO22X1_LVT U1928 ( .A1(\regs[22][27] ), .A2(n996), .A3(\regs[29][27] ), .A4(
        n973), .Y(n2725) );
  AO22X1_LVT U1929 ( .A1(\regs[2][27] ), .A2(n1014), .A3(\regs[8][27] ), .A4(
        n981), .Y(n2724) );
  AO22X1_LVT U1930 ( .A1(\regs[19][27] ), .A2(n1017), .A3(\regs[12][27] ), 
        .A4(n983), .Y(n2723) );
  NOR4X1_LVT U1931 ( .A1(n2726), .A2(n2725), .A3(n2724), .A4(n2723), .Y(n2733)
         );
  AO22X1_LVT U1932 ( .A1(\regs[31][27] ), .A2(n3481), .A3(\regs[7][27] ), .A4(
        n985), .Y(n2731) );
  AO22X1_LVT U1933 ( .A1(\regs[17][27] ), .A2(n990), .A3(\regs[30][27] ), .A4(
        n975), .Y(n2730) );
  AO22X1_LVT U1934 ( .A1(\regs[9][27] ), .A2(n967), .A3(\regs[26][27] ), .A4(
        n1002), .Y(n2729) );
  AO22X1_LVT U1935 ( .A1(\regs[3][27] ), .A2(n965), .A3(\regs[18][27] ), .A4(
        n995), .Y(n2728) );
  NOR4X1_LVT U1936 ( .A1(n2731), .A2(n2730), .A3(n2729), .A4(n2728), .Y(n2732)
         );
  NAND3X0_LVT U1937 ( .A1(n2734), .A2(n2733), .A3(n2732), .Y(n2735) );
  OR3X1_LVT U1938 ( .A1(n2737), .A2(n2736), .A3(n2735), .Y(n2738) );
  AO22X1_LVT U1939 ( .A1(wdata[27]), .A2(n960), .A3(n963), .A4(n2738), .Y(
        rdata1[27]) );
  AO22X1_LVT U1941 ( .A1(\regs[22][28] ), .A2(n996), .A3(\regs[8][28] ), .A4(
        n981), .Y(n2768) );
  AO22X1_LVT U1942 ( .A1(\regs[31][28] ), .A2(n3481), .A3(\regs[14][28] ), 
        .A4(n997), .Y(n2740) );
  INVX1_LVT U1943 ( .A(n2740), .Y(n2745) );
  AO22X1_LVT U1944 ( .A1(\regs[19][28] ), .A2(n1017), .A3(\regs[18][28] ), 
        .A4(n995), .Y(n2742) );
  INVX1_LVT U1945 ( .A(n2742), .Y(n2744) );
  NAND2X0_LVT U1946 ( .A1(\regs[11][28] ), .A2(n1022), .Y(n2743) );
  NAND3X0_LVT U1947 ( .A1(n2745), .A2(n2744), .A3(n2743), .Y(n2767) );
  AO22X1_LVT U1948 ( .A1(\regs[24][28] ), .A2(n1005), .A3(\regs[30][28] ), 
        .A4(n975), .Y(n2753) );
  AO22X1_LVT U1949 ( .A1(\regs[17][28] ), .A2(n990), .A3(\regs[3][28] ), .A4(
        n965), .Y(n2752) );
  AO22X1_LVT U1950 ( .A1(\regs[25][28] ), .A2(n979), .A3(\regs[26][28] ), .A4(
        n1002), .Y(n2751) );
  AO22X1_LVT U1951 ( .A1(\regs[7][28] ), .A2(n985), .A3(\regs[12][28] ), .A4(
        n983), .Y(n2750) );
  NOR4X1_LVT U1952 ( .A1(n2753), .A2(n2752), .A3(n2751), .A4(n2750), .Y(n2765)
         );
  AO22X1_LVT U1953 ( .A1(\regs[28][28] ), .A2(n986), .A3(\regs[21][28] ), .A4(
        n3475), .Y(n2758) );
  AO22X1_LVT U1954 ( .A1(\regs[10][28] ), .A2(n972), .A3(\regs[15][28] ), .A4(
        n1015), .Y(n2757) );
  AO22X1_LVT U1955 ( .A1(\regs[4][28] ), .A2(n1012), .A3(\regs[23][28] ), .A4(
        n968), .Y(n2756) );
  AO22X1_LVT U1956 ( .A1(\regs[29][28] ), .A2(n973), .A3(\regs[9][28] ), .A4(
        n967), .Y(n2755) );
  NOR4X1_LVT U1957 ( .A1(n2758), .A2(n2757), .A3(n2756), .A4(n2755), .Y(n2764)
         );
  AO22X1_LVT U1958 ( .A1(\regs[6][28] ), .A2(n1020), .A3(\regs[1][28] ), .A4(
        n998), .Y(n2762) );
  AO22X1_LVT U1959 ( .A1(\regs[16][28] ), .A2(n1003), .A3(\regs[5][28] ), .A4(
        n987), .Y(n2761) );
  AO22X1_LVT U1960 ( .A1(\regs[20][28] ), .A2(n1001), .A3(\regs[27][28] ), 
        .A4(n982), .Y(n2760) );
  AO22X1_LVT U1961 ( .A1(\regs[2][28] ), .A2(n1014), .A3(\regs[13][28] ), .A4(
        n1025), .Y(n2759) );
  NOR4X1_LVT U1962 ( .A1(n2762), .A2(n2761), .A3(n2760), .A4(n2759), .Y(n2763)
         );
  NAND3X0_LVT U1963 ( .A1(n2765), .A2(n2764), .A3(n2763), .Y(n2766) );
  OR3X1_LVT U1964 ( .A1(n2768), .A2(n2767), .A3(n2766), .Y(n2769) );
  AO22X1_LVT U1965 ( .A1(wdata[28]), .A2(n960), .A3(n963), .A4(n2769), .Y(
        rdata1[28]) );
  AO22X1_LVT U1967 ( .A1(\regs[26][29] ), .A2(n1002), .A3(\regs[16][29] ), 
        .A4(n1003), .Y(n2802) );
  AO22X1_LVT U1968 ( .A1(\regs[30][29] ), .A2(n975), .A3(\regs[23][29] ), .A4(
        n968), .Y(n2771) );
  INVX1_LVT U1969 ( .A(n2771), .Y(n2776) );
  AO22X1_LVT U1970 ( .A1(\regs[1][29] ), .A2(n998), .A3(\regs[31][29] ), .A4(
        n3481), .Y(n2773) );
  INVX1_LVT U1971 ( .A(n2773), .Y(n2775) );
  NAND2X0_LVT U1972 ( .A1(\regs[22][29] ), .A2(n996), .Y(n2774) );
  NAND3X0_LVT U1973 ( .A1(n2776), .A2(n2775), .A3(n2774), .Y(n2801) );
  AO22X1_LVT U1974 ( .A1(\regs[6][29] ), .A2(n1020), .A3(\regs[2][29] ), .A4(
        n1014), .Y(n2782) );
  AO22X1_LVT U1975 ( .A1(\regs[20][29] ), .A2(n1001), .A3(\regs[9][29] ), .A4(
        n967), .Y(n2781) );
  AO22X1_LVT U1976 ( .A1(\regs[8][29] ), .A2(n981), .A3(\regs[13][29] ), .A4(
        n1025), .Y(n2780) );
  AO22X1_LVT U1978 ( .A1(\regs[17][29] ), .A2(n990), .A3(\regs[15][29] ), .A4(
        n1015), .Y(n2779) );
  NOR4X1_LVT U1979 ( .A1(n2782), .A2(n2781), .A3(n2780), .A4(n2779), .Y(n2799)
         );
  AO22X1_LVT U1980 ( .A1(\regs[25][29] ), .A2(n979), .A3(\regs[18][29] ), .A4(
        n995), .Y(n2790) );
  AO22X1_LVT U1981 ( .A1(\regs[3][29] ), .A2(n965), .A3(\regs[27][29] ), .A4(
        n982), .Y(n2789) );
  AO22X1_LVT U1982 ( .A1(\regs[11][29] ), .A2(n1022), .A3(\regs[7][29] ), .A4(
        n985), .Y(n2788) );
  AO22X1_LVT U1983 ( .A1(\regs[14][29] ), .A2(n997), .A3(\regs[10][29] ), .A4(
        n972), .Y(n2787) );
  NOR4X1_LVT U1984 ( .A1(n2790), .A2(n2789), .A3(n2788), .A4(n2787), .Y(n2798)
         );
  AO22X1_LVT U1985 ( .A1(\regs[21][29] ), .A2(n3475), .A3(\regs[28][29] ), 
        .A4(n986), .Y(n2796) );
  AO22X1_LVT U1986 ( .A1(\regs[19][29] ), .A2(n1017), .A3(\regs[12][29] ), 
        .A4(n983), .Y(n2795) );
  AO22X1_LVT U1987 ( .A1(\regs[5][29] ), .A2(n987), .A3(\regs[29][29] ), .A4(
        n973), .Y(n2794) );
  AO22X1_LVT U1988 ( .A1(\regs[4][29] ), .A2(n1012), .A3(\regs[24][29] ), .A4(
        n1005), .Y(n2793) );
  NOR4X1_LVT U1989 ( .A1(n2796), .A2(n2795), .A3(n2794), .A4(n2793), .Y(n2797)
         );
  NAND3X0_LVT U1990 ( .A1(n2799), .A2(n2798), .A3(n2797), .Y(n2800) );
  OR3X1_LVT U1991 ( .A1(n2802), .A2(n2801), .A3(n2800), .Y(n2803) );
  AO22X1_LVT U1992 ( .A1(wdata[29]), .A2(n960), .A3(n963), .A4(n2803), .Y(
        rdata1[29]) );
  AO22X1_LVT U1996 ( .A1(\regs[6][30] ), .A2(n1020), .A3(\regs[4][30] ), .A4(
        n1012), .Y(n2846) );
  AO22X1_LVT U1997 ( .A1(\regs[8][30] ), .A2(n981), .A3(\regs[30][30] ), .A4(
        n975), .Y(n2809) );
  INVX1_LVT U1998 ( .A(n2809), .Y(n2815) );
  AO22X1_LVT U1999 ( .A1(\regs[12][30] ), .A2(n983), .A3(\regs[5][30] ), .A4(
        n987), .Y(n2811) );
  INVX1_LVT U2000 ( .A(n2811), .Y(n2814) );
  NAND2X0_LVT U2001 ( .A1(\regs[15][30] ), .A2(n1015), .Y(n2813) );
  NAND3X0_LVT U2002 ( .A1(n2815), .A2(n2814), .A3(n2813), .Y(n2845) );
  AO22X1_LVT U2003 ( .A1(\regs[10][30] ), .A2(n972), .A3(\regs[28][30] ), .A4(
        n986), .Y(n2822) );
  AO22X1_LVT U2004 ( .A1(\regs[26][30] ), .A2(n1002), .A3(\regs[18][30] ), 
        .A4(n995), .Y(n2821) );
  AO22X1_LVT U2005 ( .A1(\regs[11][30] ), .A2(n1022), .A3(\regs[23][30] ), 
        .A4(n968), .Y(n2820) );
  AO22X1_LVT U2007 ( .A1(\regs[21][30] ), .A2(n3475), .A3(\regs[19][30] ), 
        .A4(n1017), .Y(n2819) );
  NOR4X1_LVT U2008 ( .A1(n2822), .A2(n2821), .A3(n2820), .A4(n2819), .Y(n2843)
         );
  AO22X1_LVT U2009 ( .A1(\regs[25][30] ), .A2(n979), .A3(\regs[14][30] ), .A4(
        n997), .Y(n2832) );
  AO22X1_LVT U2010 ( .A1(\regs[7][30] ), .A2(n985), .A3(\regs[17][30] ), .A4(
        n990), .Y(n2831) );
  AO22X1_LVT U2011 ( .A1(\regs[2][30] ), .A2(n1014), .A3(\regs[27][30] ), .A4(
        n982), .Y(n2830) );
  AO22X1_LVT U2012 ( .A1(\regs[20][30] ), .A2(n1001), .A3(\regs[31][30] ), 
        .A4(n3481), .Y(n2829) );
  NOR4X1_LVT U2013 ( .A1(n2832), .A2(n2831), .A3(n2830), .A4(n2829), .Y(n2842)
         );
  AO22X1_LVT U2014 ( .A1(\regs[22][30] ), .A2(n996), .A3(\regs[24][30] ), .A4(
        n1005), .Y(n2840) );
  AO22X1_LVT U2015 ( .A1(\regs[9][30] ), .A2(n967), .A3(\regs[3][30] ), .A4(
        n965), .Y(n2839) );
  AO22X1_LVT U2016 ( .A1(\regs[13][30] ), .A2(n1025), .A3(\regs[16][30] ), 
        .A4(n1003), .Y(n2838) );
  AO22X1_LVT U2017 ( .A1(\regs[29][30] ), .A2(n973), .A3(\regs[1][30] ), .A4(
        n998), .Y(n2837) );
  NOR4X1_LVT U2018 ( .A1(n2840), .A2(n2839), .A3(n2838), .A4(n2837), .Y(n2841)
         );
  NAND3X0_LVT U2019 ( .A1(n2843), .A2(n2842), .A3(n2841), .Y(n2844) );
  OR3X1_LVT U2020 ( .A1(n2846), .A2(n2845), .A3(n2844), .Y(n2847) );
  AO22X1_LVT U2021 ( .A1(wdata[30]), .A2(n960), .A3(n963), .A4(n2847), .Y(
        rdata1[30]) );
  AO22X1_LVT U2023 ( .A1(\regs[16][31] ), .A2(n1003), .A3(\regs[29][31] ), 
        .A4(n973), .Y(n2901) );
  AO22X1_LVT U2024 ( .A1(\regs[8][31] ), .A2(n981), .A3(\regs[2][31] ), .A4(
        n1014), .Y(n2852) );
  INVX1_LVT U2025 ( .A(n2852), .Y(n2859) );
  AO22X1_LVT U2026 ( .A1(\regs[21][31] ), .A2(n3475), .A3(\regs[20][31] ), 
        .A4(n1001), .Y(n2855) );
  INVX1_LVT U2027 ( .A(n2855), .Y(n2858) );
  NAND2X0_LVT U2028 ( .A1(\regs[23][31] ), .A2(n968), .Y(n2857) );
  NAND3X0_LVT U2029 ( .A1(n2859), .A2(n2858), .A3(n2857), .Y(n2900) );
  AO22X1_LVT U2030 ( .A1(\regs[10][31] ), .A2(n972), .A3(\regs[1][31] ), .A4(
        n998), .Y(n2871) );
  AO22X1_LVT U2031 ( .A1(\regs[28][31] ), .A2(n986), .A3(\regs[30][31] ), .A4(
        n975), .Y(n2870) );
  AO22X1_LVT U2032 ( .A1(\regs[17][31] ), .A2(n990), .A3(\regs[22][31] ), .A4(
        n996), .Y(n2869) );
  AO22X1_LVT U2033 ( .A1(\regs[4][31] ), .A2(n1012), .A3(\regs[25][31] ), .A4(
        n979), .Y(n2868) );
  NOR4X1_LVT U2034 ( .A1(n2871), .A2(n2870), .A3(n2869), .A4(n2868), .Y(n2898)
         );
  AO22X1_LVT U2035 ( .A1(\regs[15][31] ), .A2(n1015), .A3(\regs[7][31] ), .A4(
        n985), .Y(n2883) );
  AO22X1_LVT U2036 ( .A1(\regs[5][31] ), .A2(n987), .A3(\regs[18][31] ), .A4(
        n995), .Y(n2882) );
  AO22X1_LVT U2037 ( .A1(\regs[13][31] ), .A2(n1025), .A3(\regs[19][31] ), 
        .A4(n1017), .Y(n2881) );
  AO22X1_LVT U2038 ( .A1(\regs[26][31] ), .A2(n1002), .A3(\regs[24][31] ), 
        .A4(n1005), .Y(n2880) );
  NOR4X1_LVT U2039 ( .A1(n2883), .A2(n2882), .A3(n2881), .A4(n2880), .Y(n2897)
         );
  AO22X1_LVT U2040 ( .A1(\regs[12][31] ), .A2(n983), .A3(\regs[11][31] ), .A4(
        n1022), .Y(n2895) );
  AO22X1_LVT U2041 ( .A1(\regs[31][31] ), .A2(n3481), .A3(\regs[27][31] ), 
        .A4(n982), .Y(n2894) );
  AO22X1_LVT U2042 ( .A1(\regs[14][31] ), .A2(n997), .A3(\regs[3][31] ), .A4(
        n965), .Y(n2893) );
  AO22X1_LVT U2043 ( .A1(\regs[6][31] ), .A2(n1020), .A3(\regs[9][31] ), .A4(
        n967), .Y(n2892) );
  NOR4X1_LVT U2044 ( .A1(n2895), .A2(n2894), .A3(n2893), .A4(n2892), .Y(n2896)
         );
  NAND3X0_LVT U2045 ( .A1(n2898), .A2(n2897), .A3(n2896), .Y(n2899) );
  OR3X1_LVT U2046 ( .A1(n2901), .A2(n2900), .A3(n2899), .Y(n2902) );
  AO22X1_LVT U2047 ( .A1(wdata[31]), .A2(n960), .A3(n963), .A4(n2902), .Y(
        rdata1[31]) );
  AND2X2_LVT U2048 ( .A1(waddr[0]), .A2(n3192), .Y(n3202) );
  AND4X1_LVT U2049 ( .A1(we), .A2(n3077), .A3(n3002), .A4(n3297), .Y(n2992) );
  AND2X1_LVT U2050 ( .A1(n2992), .A2(n3298), .Y(n2955) );
  AO22X1_LVT U2056 ( .A1(n3443), .A2(n3486), .A3(n3442), .A4(\regs[1][31] ), 
        .Y(n2530) );
  AO22X1_LVT U2057 ( .A1(n3443), .A2(wdata[30]), .A3(n3442), .A4(\regs[1][30] ), .Y(n2529) );
  AO22X1_LVT U2058 ( .A1(n3443), .A2(n3501), .A3(n3442), .A4(\regs[1][29] ), 
        .Y(n2528) );
  AO22X1_LVT U2059 ( .A1(n3443), .A2(n3500), .A3(n3442), .A4(\regs[1][28] ), 
        .Y(n2527) );
  AO22X1_LVT U2060 ( .A1(n3443), .A2(wdata[27]), .A3(n3442), .A4(\regs[1][27] ), .Y(n2526) );
  AO22X1_LVT U2061 ( .A1(n3443), .A2(n3503), .A3(n3442), .A4(\regs[1][26] ), 
        .Y(n2525) );
  AO22X1_LVT U2062 ( .A1(n3443), .A2(wdata[25]), .A3(n3442), .A4(\regs[1][25] ), .Y(n2524) );
  AO22X1_LVT U2064 ( .A1(n3447), .A2(n3493), .A3(n3446), .A4(\regs[1][24] ), 
        .Y(n2523) );
  AO22X1_LVT U2065 ( .A1(n3447), .A2(n3497), .A3(n3446), .A4(\regs[1][23] ), 
        .Y(n2522) );
  AO22X1_LVT U2066 ( .A1(n3447), .A2(n3494), .A3(n3446), .A4(\regs[1][22] ), 
        .Y(n2521) );
  AO22X1_LVT U2067 ( .A1(n3447), .A2(wdata[21]), .A3(n3446), .A4(\regs[1][21] ), .Y(n2520) );
  AO22X1_LVT U2068 ( .A1(n3447), .A2(n3483), .A3(n3446), .A4(\regs[1][20] ), 
        .Y(n2519) );
  AO22X1_LVT U2069 ( .A1(n3447), .A2(n3496), .A3(n3446), .A4(\regs[1][19] ), 
        .Y(n2518) );
  AO22X1_LVT U2070 ( .A1(n3447), .A2(n3491), .A3(n3446), .A4(\regs[1][18] ), 
        .Y(n2517) );
  AO22X1_LVT U2071 ( .A1(n3447), .A2(wdata[17]), .A3(n3446), .A4(\regs[1][17] ), .Y(n2516) );
  AO22X1_LVT U2073 ( .A1(n3443), .A2(wdata[16]), .A3(n3442), .A4(\regs[1][16] ), .Y(n2515) );
  AO22X1_LVT U2074 ( .A1(n3443), .A2(n3495), .A3(n3442), .A4(\regs[1][15] ), 
        .Y(n2514) );
  AO22X1_LVT U2075 ( .A1(n3443), .A2(n3498), .A3(n3442), .A4(\regs[1][14] ), 
        .Y(n2513) );
  AO22X1_LVT U2076 ( .A1(n3443), .A2(n3502), .A3(n3442), .A4(\regs[1][13] ), 
        .Y(n2512) );
  AO22X1_LVT U2077 ( .A1(n3443), .A2(wdata[12]), .A3(n3442), .A4(\regs[1][12] ), .Y(n2511) );
  AO22X1_LVT U2078 ( .A1(n3443), .A2(wdata[11]), .A3(n3442), .A4(\regs[1][11] ), .Y(n2510) );
  AO22X1_LVT U2079 ( .A1(n3443), .A2(n3499), .A3(n3442), .A4(\regs[1][10] ), 
        .Y(n2509) );
  AO22X1_LVT U2080 ( .A1(n3443), .A2(wdata[9]), .A3(n3442), .A4(\regs[1][9] ), 
        .Y(n2508) );
  AO22X1_LVT U2082 ( .A1(n3445), .A2(wdata[8]), .A3(n3444), .A4(\regs[1][8] ), 
        .Y(n2507) );
  AO22X1_LVT U2083 ( .A1(n3445), .A2(wdata[7]), .A3(n3444), .A4(\regs[1][7] ), 
        .Y(n2506) );
  AO22X1_LVT U2084 ( .A1(n3445), .A2(wdata[6]), .A3(n3444), .A4(\regs[1][6] ), 
        .Y(n2505) );
  AO22X1_LVT U2085 ( .A1(n3445), .A2(wdata[5]), .A3(n3444), .A4(\regs[1][5] ), 
        .Y(n2504) );
  AO22X1_LVT U2086 ( .A1(n3445), .A2(wdata[4]), .A3(n3444), .A4(\regs[1][4] ), 
        .Y(n2503) );
  AO22X1_LVT U2087 ( .A1(n3445), .A2(wdata[3]), .A3(n3444), .A4(\regs[1][3] ), 
        .Y(n2502) );
  AO22X1_LVT U2088 ( .A1(n3445), .A2(wdata[2]), .A3(n3444), .A4(\regs[1][2] ), 
        .Y(n2501) );
  AO22X1_LVT U2090 ( .A1(n3445), .A2(wdata[1]), .A3(n3444), .A4(\regs[1][1] ), 
        .Y(n2500) );
  AO22X1_LVT U2091 ( .A1(n3445), .A2(wdata[0]), .A3(n3444), .A4(\regs[1][0] ), 
        .Y(n2499) );
  AND2X2_LVT U2092 ( .A1(waddr[1]), .A2(n3191), .Y(n3212) );
  AO22X1_LVT U2098 ( .A1(n3437), .A2(n3486), .A3(n3436), .A4(\regs[2][31] ), 
        .Y(n2498) );
  AO22X1_LVT U2099 ( .A1(n3437), .A2(wdata[30]), .A3(n3436), .A4(\regs[2][30] ), .Y(n2497) );
  AO22X1_LVT U2100 ( .A1(n3437), .A2(n3501), .A3(n3436), .A4(\regs[2][29] ), 
        .Y(n2496) );
  AO22X1_LVT U2101 ( .A1(n3437), .A2(n3500), .A3(n3436), .A4(\regs[2][28] ), 
        .Y(n2495) );
  AO22X1_LVT U2102 ( .A1(n3437), .A2(wdata[27]), .A3(n3436), .A4(\regs[2][27] ), .Y(n2494) );
  AO22X1_LVT U2103 ( .A1(n3437), .A2(wdata[26]), .A3(n3436), .A4(\regs[2][26] ), .Y(n2493) );
  AO22X1_LVT U2104 ( .A1(n3437), .A2(wdata[25]), .A3(n3436), .A4(\regs[2][25] ), .Y(n2492) );
  AO22X1_LVT U2106 ( .A1(n3441), .A2(n3493), .A3(n3440), .A4(\regs[2][24] ), 
        .Y(n2491) );
  AO22X1_LVT U2107 ( .A1(n3441), .A2(n3497), .A3(n3440), .A4(\regs[2][23] ), 
        .Y(n2490) );
  AO22X1_LVT U2108 ( .A1(n3441), .A2(n3494), .A3(n3440), .A4(\regs[2][22] ), 
        .Y(n2489) );
  AO22X1_LVT U2109 ( .A1(n3441), .A2(wdata[21]), .A3(n3440), .A4(\regs[2][21] ), .Y(n2488) );
  AO22X1_LVT U2110 ( .A1(n3441), .A2(n3483), .A3(n3440), .A4(\regs[2][20] ), 
        .Y(n2487) );
  AO22X1_LVT U2111 ( .A1(n3441), .A2(n3496), .A3(n3440), .A4(\regs[2][19] ), 
        .Y(n2486) );
  AO22X1_LVT U2112 ( .A1(n3441), .A2(n3491), .A3(n3440), .A4(\regs[2][18] ), 
        .Y(n2485) );
  AO22X1_LVT U2113 ( .A1(n3441), .A2(wdata[17]), .A3(n3440), .A4(\regs[2][17] ), .Y(n2484) );
  AO22X1_LVT U2115 ( .A1(n3437), .A2(wdata[16]), .A3(n3436), .A4(\regs[2][16] ), .Y(n2483) );
  AO22X1_LVT U2116 ( .A1(n3441), .A2(n3495), .A3(n3440), .A4(\regs[2][15] ), 
        .Y(n2482) );
  AO22X1_LVT U2117 ( .A1(n3441), .A2(n3498), .A3(n3440), .A4(\regs[2][14] ), 
        .Y(n2481) );
  AO22X1_LVT U2118 ( .A1(n3437), .A2(n3502), .A3(n3436), .A4(\regs[2][13] ), 
        .Y(n2480) );
  AO22X1_LVT U2119 ( .A1(n3437), .A2(wdata[12]), .A3(n3436), .A4(\regs[2][12] ), .Y(n2479) );
  AO22X1_LVT U2120 ( .A1(n3437), .A2(wdata[11]), .A3(n3436), .A4(\regs[2][11] ), .Y(n2478) );
  AO22X1_LVT U2121 ( .A1(n3437), .A2(n3499), .A3(n3436), .A4(\regs[2][10] ), 
        .Y(n2477) );
  AO22X1_LVT U2122 ( .A1(n3437), .A2(wdata[9]), .A3(n3436), .A4(\regs[2][9] ), 
        .Y(n2476) );
  AO22X1_LVT U2124 ( .A1(n3439), .A2(wdata[8]), .A3(n3438), .A4(\regs[2][8] ), 
        .Y(n2475) );
  AO22X1_LVT U2125 ( .A1(n3439), .A2(wdata[7]), .A3(n3438), .A4(\regs[2][7] ), 
        .Y(n2474) );
  AO22X1_LVT U2126 ( .A1(n3439), .A2(wdata[6]), .A3(n3438), .A4(\regs[2][6] ), 
        .Y(n2473) );
  AO22X1_LVT U2127 ( .A1(n3439), .A2(wdata[5]), .A3(n3438), .A4(\regs[2][5] ), 
        .Y(n2472) );
  AO22X1_LVT U2128 ( .A1(n3439), .A2(wdata[4]), .A3(n3438), .A4(\regs[2][4] ), 
        .Y(n2471) );
  AO22X1_LVT U2129 ( .A1(n3439), .A2(wdata[3]), .A3(n3438), .A4(\regs[2][3] ), 
        .Y(n2470) );
  AO22X1_LVT U2130 ( .A1(n3439), .A2(wdata[2]), .A3(n3438), .A4(\regs[2][2] ), 
        .Y(n2469) );
  AO22X1_LVT U2132 ( .A1(n3439), .A2(wdata[1]), .A3(n3438), .A4(\regs[2][1] ), 
        .Y(n2468) );
  AO22X1_LVT U2133 ( .A1(n3439), .A2(wdata[0]), .A3(n3438), .A4(\regs[2][0] ), 
        .Y(n2467) );
  NAND2X0_LVT U2135 ( .A1(n2955), .A2(n3255), .Y(n2956) );
  AO22X1_LVT U2141 ( .A1(n3435), .A2(n3486), .A3(n3434), .A4(\regs[3][31] ), 
        .Y(n2466) );
  AO22X1_LVT U2143 ( .A1(n3435), .A2(wdata[30]), .A3(n3434), .A4(\regs[3][30] ), .Y(n2465) );
  AO22X1_LVT U2145 ( .A1(n3435), .A2(n3501), .A3(n3434), .A4(\regs[3][29] ), 
        .Y(n2464) );
  AO22X1_LVT U2147 ( .A1(n3435), .A2(n3500), .A3(n3434), .A4(\regs[3][28] ), 
        .Y(n2463) );
  AO22X1_LVT U2149 ( .A1(n3435), .A2(wdata[27]), .A3(n3434), .A4(\regs[3][27] ), .Y(n2462) );
  AO22X1_LVT U2151 ( .A1(n3435), .A2(n3503), .A3(n3434), .A4(\regs[3][26] ), 
        .Y(n2461) );
  AO22X1_LVT U2153 ( .A1(n3435), .A2(wdata[25]), .A3(n3434), .A4(\regs[3][25] ), .Y(n2460) );
  AO22X1_LVT U2156 ( .A1(n3433), .A2(n3493), .A3(n3432), .A4(\regs[3][24] ), 
        .Y(n2459) );
  AO22X1_LVT U2158 ( .A1(n3433), .A2(n3497), .A3(n3432), .A4(\regs[3][23] ), 
        .Y(n2458) );
  AO22X1_LVT U2160 ( .A1(n3433), .A2(n3494), .A3(n3432), .A4(\regs[3][22] ), 
        .Y(n2457) );
  AO22X1_LVT U2162 ( .A1(n3433), .A2(wdata[21]), .A3(n3432), .A4(\regs[3][21] ), .Y(n2456) );
  AO22X1_LVT U2164 ( .A1(n3433), .A2(n3483), .A3(n3432), .A4(\regs[3][20] ), 
        .Y(n2455) );
  AO22X1_LVT U2166 ( .A1(n3433), .A2(n3496), .A3(n3432), .A4(\regs[3][19] ), 
        .Y(n2454) );
  AO22X1_LVT U2168 ( .A1(n3433), .A2(n3491), .A3(n3432), .A4(\regs[3][18] ), 
        .Y(n2453) );
  AO22X1_LVT U2170 ( .A1(n3433), .A2(wdata[17]), .A3(n3432), .A4(\regs[3][17] ), .Y(n2452) );
  AO22X1_LVT U2173 ( .A1(n3435), .A2(wdata[16]), .A3(n3434), .A4(\regs[3][16] ), .Y(n2451) );
  AO22X1_LVT U2175 ( .A1(n3435), .A2(n3495), .A3(n3434), .A4(\regs[3][15] ), 
        .Y(n2450) );
  AO22X1_LVT U2177 ( .A1(n3435), .A2(n3498), .A3(n3434), .A4(\regs[3][14] ), 
        .Y(n2449) );
  AO22X1_LVT U2179 ( .A1(n3435), .A2(n3502), .A3(n3434), .A4(\regs[3][13] ), 
        .Y(n2448) );
  AO22X1_LVT U2181 ( .A1(n3435), .A2(wdata[12]), .A3(n3434), .A4(\regs[3][12] ), .Y(n2447) );
  AO22X1_LVT U2183 ( .A1(n3435), .A2(wdata[11]), .A3(n3434), .A4(\regs[3][11] ), .Y(n2446) );
  AO22X1_LVT U2185 ( .A1(n3435), .A2(n3499), .A3(n3434), .A4(\regs[3][10] ), 
        .Y(n2445) );
  AO22X1_LVT U2187 ( .A1(n3435), .A2(wdata[9]), .A3(n3434), .A4(\regs[3][9] ), 
        .Y(n2444) );
  AO22X1_LVT U2190 ( .A1(n3433), .A2(wdata[8]), .A3(n3432), .A4(\regs[3][8] ), 
        .Y(n2443) );
  AO22X1_LVT U2192 ( .A1(n3433), .A2(wdata[7]), .A3(n3432), .A4(\regs[3][7] ), 
        .Y(n2442) );
  AO22X1_LVT U2194 ( .A1(n3433), .A2(wdata[6]), .A3(n3432), .A4(\regs[3][6] ), 
        .Y(n2441) );
  AO22X1_LVT U2196 ( .A1(n3433), .A2(wdata[5]), .A3(n3432), .A4(\regs[3][5] ), 
        .Y(n2440) );
  AO22X1_LVT U2198 ( .A1(n3433), .A2(wdata[4]), .A3(n3432), .A4(\regs[3][4] ), 
        .Y(n2439) );
  AO22X1_LVT U2200 ( .A1(n3433), .A2(wdata[3]), .A3(n3432), .A4(\regs[3][3] ), 
        .Y(n2438) );
  AO22X1_LVT U2202 ( .A1(n3433), .A2(wdata[2]), .A3(n3432), .A4(\regs[3][2] ), 
        .Y(n2437) );
  AO22X1_LVT U2205 ( .A1(n3433), .A2(wdata[1]), .A3(n3432), .A4(\regs[3][1] ), 
        .Y(n2436) );
  AO22X1_LVT U2207 ( .A1(n3433), .A2(wdata[0]), .A3(n3432), .A4(\regs[3][0] ), 
        .Y(n2435) );
  NAND4X0_LVT U2208 ( .A1(n3470), .A2(n2992), .A3(n3192), .A4(n3191), .Y(n2965) );
  AO22X1_LVT U2213 ( .A1(n3316), .A2(n3486), .A3(n3315), .A4(\regs[4][31] ), 
        .Y(n2434) );
  AO22X1_LVT U2214 ( .A1(n3316), .A2(wdata[30]), .A3(n3315), .A4(\regs[4][30] ), .Y(n2433) );
  AO22X1_LVT U2215 ( .A1(n3316), .A2(n3501), .A3(n3315), .A4(\regs[4][29] ), 
        .Y(n2432) );
  AO22X1_LVT U2216 ( .A1(n3316), .A2(n3500), .A3(n3315), .A4(\regs[4][28] ), 
        .Y(n2431) );
  AO22X1_LVT U2217 ( .A1(n3316), .A2(wdata[27]), .A3(n3315), .A4(\regs[4][27] ), .Y(n2430) );
  AO22X1_LVT U2218 ( .A1(n3316), .A2(n3503), .A3(n3315), .A4(\regs[4][26] ), 
        .Y(n2429) );
  AO22X1_LVT U2219 ( .A1(n3316), .A2(wdata[25]), .A3(n3315), .A4(\regs[4][25] ), .Y(n2428) );
  AO22X1_LVT U2221 ( .A1(n3318), .A2(n3493), .A3(n3317), .A4(\regs[4][24] ), 
        .Y(n2427) );
  AO22X1_LVT U2222 ( .A1(n3316), .A2(n3497), .A3(n3315), .A4(\regs[4][23] ), 
        .Y(n2426) );
  AO22X1_LVT U2223 ( .A1(n3318), .A2(n3494), .A3(n3317), .A4(\regs[4][22] ), 
        .Y(n2425) );
  AO22X1_LVT U2224 ( .A1(n3316), .A2(wdata[21]), .A3(n3315), .A4(\regs[4][21] ), .Y(n2424) );
  AO22X1_LVT U2225 ( .A1(n3318), .A2(n3483), .A3(n3317), .A4(\regs[4][20] ), 
        .Y(n2423) );
  AO22X1_LVT U2226 ( .A1(n3316), .A2(n3496), .A3(n3315), .A4(\regs[4][19] ), 
        .Y(n2422) );
  AO22X1_LVT U2227 ( .A1(n3318), .A2(n3491), .A3(n3317), .A4(\regs[4][18] ), 
        .Y(n2421) );
  AO22X1_LVT U2228 ( .A1(n3316), .A2(wdata[17]), .A3(n3315), .A4(\regs[4][17] ), .Y(n2420) );
  AO22X1_LVT U2230 ( .A1(n3316), .A2(wdata[16]), .A3(n3315), .A4(\regs[4][16] ), .Y(n2419) );
  AO22X1_LVT U2231 ( .A1(n3316), .A2(n3495), .A3(n3315), .A4(\regs[4][15] ), 
        .Y(n2418) );
  AO22X1_LVT U2232 ( .A1(n3316), .A2(n3498), .A3(n3315), .A4(\regs[4][14] ), 
        .Y(n2417) );
  AO22X1_LVT U2233 ( .A1(n3316), .A2(n3502), .A3(n3315), .A4(\regs[4][13] ), 
        .Y(n2416) );
  AO22X1_LVT U2234 ( .A1(n3316), .A2(wdata[12]), .A3(n3315), .A4(\regs[4][12] ), .Y(n2415) );
  AO22X1_LVT U2235 ( .A1(n3316), .A2(wdata[11]), .A3(n3315), .A4(\regs[4][11] ), .Y(n2414) );
  AO22X1_LVT U2236 ( .A1(n3316), .A2(n3499), .A3(n3315), .A4(\regs[4][10] ), 
        .Y(n2413) );
  AO22X1_LVT U2237 ( .A1(n3316), .A2(wdata[9]), .A3(n3315), .A4(\regs[4][9] ), 
        .Y(n2412) );
  AO22X1_LVT U2239 ( .A1(n3318), .A2(wdata[8]), .A3(n3317), .A4(\regs[4][8] ), 
        .Y(n2411) );
  AO22X1_LVT U2240 ( .A1(n3318), .A2(wdata[7]), .A3(n3317), .A4(\regs[4][7] ), 
        .Y(n2410) );
  AO22X1_LVT U2241 ( .A1(n3318), .A2(wdata[6]), .A3(n3317), .A4(\regs[4][6] ), 
        .Y(n2409) );
  AO22X1_LVT U2242 ( .A1(n3318), .A2(wdata[5]), .A3(n3317), .A4(\regs[4][5] ), 
        .Y(n2408) );
  AO22X1_LVT U2243 ( .A1(n3318), .A2(wdata[4]), .A3(n3317), .A4(\regs[4][4] ), 
        .Y(n2407) );
  AO22X1_LVT U2244 ( .A1(n3318), .A2(wdata[3]), .A3(n3317), .A4(\regs[4][3] ), 
        .Y(n2406) );
  AO22X1_LVT U2245 ( .A1(n3318), .A2(wdata[2]), .A3(n3317), .A4(\regs[4][2] ), 
        .Y(n2405) );
  AO22X1_LVT U2247 ( .A1(n3318), .A2(wdata[1]), .A3(n3317), .A4(\regs[4][1] ), 
        .Y(n2404) );
  AO22X1_LVT U2248 ( .A1(n3318), .A2(wdata[0]), .A3(n3317), .A4(\regs[4][0] ), 
        .Y(n2403) );
  AO22X1_LVT U2254 ( .A1(n3374), .A2(n3486), .A3(n3373), .A4(\regs[5][31] ), 
        .Y(n2402) );
  AO22X1_LVT U2255 ( .A1(n3374), .A2(wdata[30]), .A3(n3373), .A4(\regs[5][30] ), .Y(n2401) );
  AO22X1_LVT U2256 ( .A1(n3374), .A2(n3501), .A3(n3373), .A4(\regs[5][29] ), 
        .Y(n2400) );
  AO22X1_LVT U2257 ( .A1(n3374), .A2(wdata[28]), .A3(n3373), .A4(\regs[5][28] ), .Y(n2399) );
  AO22X1_LVT U2258 ( .A1(n3374), .A2(wdata[27]), .A3(n3373), .A4(\regs[5][27] ), .Y(n2398) );
  AO22X1_LVT U2259 ( .A1(n3374), .A2(n3503), .A3(n3373), .A4(\regs[5][26] ), 
        .Y(n2397) );
  AO22X1_LVT U2260 ( .A1(n3374), .A2(wdata[25]), .A3(n3373), .A4(\regs[5][25] ), .Y(n2396) );
  AO22X1_LVT U2262 ( .A1(n3378), .A2(n3493), .A3(n3377), .A4(\regs[5][24] ), 
        .Y(n2395) );
  AO22X1_LVT U2263 ( .A1(n3378), .A2(n3497), .A3(n3377), .A4(\regs[5][23] ), 
        .Y(n2394) );
  AO22X1_LVT U2264 ( .A1(n3378), .A2(n3494), .A3(n3377), .A4(\regs[5][22] ), 
        .Y(n2393) );
  AO22X1_LVT U2265 ( .A1(n3378), .A2(wdata[21]), .A3(n3377), .A4(\regs[5][21] ), .Y(n2392) );
  AO22X1_LVT U2266 ( .A1(n3378), .A2(n3483), .A3(n3377), .A4(\regs[5][20] ), 
        .Y(n2391) );
  AO22X1_LVT U2267 ( .A1(n3378), .A2(wdata[19]), .A3(n3377), .A4(\regs[5][19] ), .Y(n2390) );
  AO22X1_LVT U2268 ( .A1(n3378), .A2(n3491), .A3(n3377), .A4(\regs[5][18] ), 
        .Y(n2389) );
  AO22X1_LVT U2269 ( .A1(n3376), .A2(wdata[17]), .A3(n3377), .A4(\regs[5][17] ), .Y(n2388) );
  AO22X1_LVT U2271 ( .A1(n3374), .A2(wdata[16]), .A3(n3373), .A4(\regs[5][16] ), .Y(n2387) );
  AO22X1_LVT U2272 ( .A1(n3374), .A2(n3495), .A3(n3373), .A4(\regs[5][15] ), 
        .Y(n2386) );
  AO22X1_LVT U2273 ( .A1(n3374), .A2(n3498), .A3(n3373), .A4(\regs[5][14] ), 
        .Y(n2385) );
  AO22X1_LVT U2274 ( .A1(n3374), .A2(n3502), .A3(n3373), .A4(\regs[5][13] ), 
        .Y(n2384) );
  AO22X1_LVT U2275 ( .A1(n3374), .A2(wdata[12]), .A3(n3373), .A4(\regs[5][12] ), .Y(n2383) );
  AO22X1_LVT U2276 ( .A1(n3374), .A2(wdata[11]), .A3(n3373), .A4(\regs[5][11] ), .Y(n2382) );
  AO22X1_LVT U2277 ( .A1(n3374), .A2(n3499), .A3(n3373), .A4(\regs[5][10] ), 
        .Y(n2381) );
  AO22X1_LVT U2278 ( .A1(n3374), .A2(wdata[9]), .A3(n3373), .A4(\regs[5][9] ), 
        .Y(n2380) );
  AO22X1_LVT U2280 ( .A1(n3376), .A2(wdata[8]), .A3(n3377), .A4(\regs[5][8] ), 
        .Y(n2379) );
  AO22X1_LVT U2281 ( .A1(n3376), .A2(wdata[7]), .A3(n3377), .A4(\regs[5][7] ), 
        .Y(n2378) );
  AO22X1_LVT U2282 ( .A1(n3376), .A2(wdata[6]), .A3(n3377), .A4(\regs[5][6] ), 
        .Y(n2377) );
  AO22X1_LVT U2283 ( .A1(n3376), .A2(wdata[5]), .A3(n3377), .A4(\regs[5][5] ), 
        .Y(n2376) );
  AO22X1_LVT U2284 ( .A1(n3376), .A2(wdata[4]), .A3(n3377), .A4(\regs[5][4] ), 
        .Y(n2375) );
  AO22X1_LVT U2285 ( .A1(n3376), .A2(wdata[3]), .A3(n3377), .A4(\regs[5][3] ), 
        .Y(n2374) );
  AO22X1_LVT U2286 ( .A1(n3376), .A2(wdata[2]), .A3(n3377), .A4(\regs[5][2] ), 
        .Y(n2373) );
  AO22X1_LVT U2288 ( .A1(n3376), .A2(wdata[1]), .A3(n3377), .A4(\regs[5][1] ), 
        .Y(n2372) );
  AO22X1_LVT U2289 ( .A1(n3376), .A2(wdata[0]), .A3(n3377), .A4(\regs[5][0] ), 
        .Y(n2371) );
  AO22X1_LVT U2295 ( .A1(n3368), .A2(n3486), .A3(n3367), .A4(\regs[6][31] ), 
        .Y(n2370) );
  AO22X1_LVT U2296 ( .A1(n3368), .A2(wdata[30]), .A3(n3367), .A4(\regs[6][30] ), .Y(n2369) );
  AO22X1_LVT U2297 ( .A1(n3368), .A2(n3501), .A3(n3367), .A4(\regs[6][29] ), 
        .Y(n2368) );
  AO22X1_LVT U2298 ( .A1(n3368), .A2(n3500), .A3(n3367), .A4(\regs[6][28] ), 
        .Y(n2367) );
  AO22X1_LVT U2299 ( .A1(n3368), .A2(wdata[27]), .A3(n3367), .A4(\regs[6][27] ), .Y(n2366) );
  AO22X1_LVT U2300 ( .A1(n3368), .A2(n3503), .A3(n3367), .A4(\regs[6][26] ), 
        .Y(n2365) );
  AO22X1_LVT U2301 ( .A1(n3368), .A2(wdata[25]), .A3(n3367), .A4(\regs[6][25] ), .Y(n2364) );
  AO22X1_LVT U2303 ( .A1(n3372), .A2(n3493), .A3(n3371), .A4(\regs[6][24] ), 
        .Y(n2363) );
  AO22X1_LVT U2304 ( .A1(n3372), .A2(n3497), .A3(n3371), .A4(\regs[6][23] ), 
        .Y(n2362) );
  AO22X1_LVT U2305 ( .A1(n3372), .A2(n3494), .A3(n3371), .A4(\regs[6][22] ), 
        .Y(n2361) );
  AO22X1_LVT U2306 ( .A1(n3372), .A2(wdata[21]), .A3(n3371), .A4(\regs[6][21] ), .Y(n2360) );
  AO22X1_LVT U2307 ( .A1(n3372), .A2(n3483), .A3(n3371), .A4(\regs[6][20] ), 
        .Y(n2359) );
  AO22X1_LVT U2308 ( .A1(n3372), .A2(n3496), .A3(n3371), .A4(\regs[6][19] ), 
        .Y(n2358) );
  AO22X1_LVT U2309 ( .A1(n3372), .A2(n3491), .A3(n3371), .A4(\regs[6][18] ), 
        .Y(n2357) );
  AO22X1_LVT U2310 ( .A1(n3372), .A2(wdata[17]), .A3(n3371), .A4(\regs[6][17] ), .Y(n2356) );
  AO22X1_LVT U2312 ( .A1(n3370), .A2(wdata[16]), .A3(n3369), .A4(\regs[6][16] ), .Y(n2355) );
  AO22X1_LVT U2313 ( .A1(n3368), .A2(n3495), .A3(n3367), .A4(\regs[6][15] ), 
        .Y(n2354) );
  AO22X1_LVT U2314 ( .A1(n3370), .A2(n3498), .A3(n3369), .A4(\regs[6][14] ), 
        .Y(n2353) );
  AO22X1_LVT U2315 ( .A1(n3370), .A2(n3502), .A3(n3369), .A4(\regs[6][13] ), 
        .Y(n2352) );
  AO22X1_LVT U2316 ( .A1(n3368), .A2(wdata[12]), .A3(n3367), .A4(\regs[6][12] ), .Y(n2351) );
  AO22X1_LVT U2317 ( .A1(n3370), .A2(wdata[11]), .A3(n3369), .A4(\regs[6][11] ), .Y(n2350) );
  AO22X1_LVT U2318 ( .A1(n3370), .A2(n3499), .A3(n3369), .A4(\regs[6][10] ), 
        .Y(n2349) );
  AO22X1_LVT U2319 ( .A1(n3370), .A2(wdata[9]), .A3(n3369), .A4(\regs[6][9] ), 
        .Y(n2348) );
  AO22X1_LVT U2321 ( .A1(n3372), .A2(wdata[8]), .A3(n3371), .A4(\regs[6][8] ), 
        .Y(n2347) );
  AO22X1_LVT U2322 ( .A1(n3370), .A2(wdata[7]), .A3(n3369), .A4(\regs[6][7] ), 
        .Y(n2346) );
  AO22X1_LVT U2323 ( .A1(n3370), .A2(wdata[6]), .A3(n3369), .A4(\regs[6][6] ), 
        .Y(n2345) );
  AO22X1_LVT U2324 ( .A1(n3372), .A2(wdata[5]), .A3(n3371), .A4(\regs[6][5] ), 
        .Y(n2344) );
  AO22X1_LVT U2325 ( .A1(n3370), .A2(wdata[4]), .A3(n3369), .A4(\regs[6][4] ), 
        .Y(n2343) );
  AO22X1_LVT U2326 ( .A1(n3372), .A2(wdata[3]), .A3(n3371), .A4(\regs[6][3] ), 
        .Y(n2342) );
  AO22X1_LVT U2327 ( .A1(n3372), .A2(wdata[2]), .A3(n3371), .A4(\regs[6][2] ), 
        .Y(n2341) );
  AO22X1_LVT U2329 ( .A1(n3372), .A2(wdata[1]), .A3(n3371), .A4(\regs[6][1] ), 
        .Y(n2340) );
  AO22X1_LVT U2330 ( .A1(n3372), .A2(wdata[0]), .A3(n3371), .A4(\regs[6][0] ), 
        .Y(n2339) );
  AO22X1_LVT U2336 ( .A1(n3364), .A2(n3486), .A3(n3363), .A4(\regs[7][31] ), 
        .Y(n2338) );
  AO22X1_LVT U2337 ( .A1(n3364), .A2(wdata[30]), .A3(n3363), .A4(\regs[7][30] ), .Y(n2337) );
  AO22X1_LVT U2338 ( .A1(n3364), .A2(n3501), .A3(n3363), .A4(\regs[7][29] ), 
        .Y(n2336) );
  AO22X1_LVT U2339 ( .A1(n3364), .A2(n3500), .A3(n3363), .A4(\regs[7][28] ), 
        .Y(n2335) );
  AO22X1_LVT U2340 ( .A1(n3364), .A2(wdata[27]), .A3(n3363), .A4(\regs[7][27] ), .Y(n2334) );
  AO22X1_LVT U2341 ( .A1(n3364), .A2(n3503), .A3(n3363), .A4(\regs[7][26] ), 
        .Y(n2333) );
  AO22X1_LVT U2342 ( .A1(n3364), .A2(wdata[25]), .A3(n3363), .A4(\regs[7][25] ), .Y(n2332) );
  AO22X1_LVT U2344 ( .A1(n3366), .A2(n3493), .A3(n3363), .A4(\regs[7][24] ), 
        .Y(n2331) );
  AO22X1_LVT U2345 ( .A1(n3366), .A2(n3497), .A3(n3363), .A4(\regs[7][23] ), 
        .Y(n2330) );
  AO22X1_LVT U2346 ( .A1(n3362), .A2(n3494), .A3(n3363), .A4(\regs[7][22] ), 
        .Y(n2329) );
  AO22X1_LVT U2347 ( .A1(n3366), .A2(wdata[21]), .A3(n3363), .A4(\regs[7][21] ), .Y(n2328) );
  AO22X1_LVT U2348 ( .A1(n3366), .A2(n3483), .A3(n3363), .A4(\regs[7][20] ), 
        .Y(n2327) );
  AO22X1_LVT U2349 ( .A1(n3366), .A2(n3496), .A3(n3363), .A4(\regs[7][19] ), 
        .Y(n2326) );
  AO22X1_LVT U2350 ( .A1(n3366), .A2(n3491), .A3(n3363), .A4(\regs[7][18] ), 
        .Y(n2325) );
  AO22X1_LVT U2351 ( .A1(n3362), .A2(wdata[17]), .A3(n3363), .A4(\regs[7][17] ), .Y(n2324) );
  AO22X1_LVT U2353 ( .A1(n3364), .A2(wdata[16]), .A3(n3363), .A4(\regs[7][16] ), .Y(n2323) );
  AO22X1_LVT U2354 ( .A1(n3364), .A2(n3495), .A3(n3363), .A4(\regs[7][15] ), 
        .Y(n2322) );
  AO22X1_LVT U2355 ( .A1(n3364), .A2(n3498), .A3(n3363), .A4(\regs[7][14] ), 
        .Y(n2321) );
  AO22X1_LVT U2356 ( .A1(n3364), .A2(n3502), .A3(n3363), .A4(\regs[7][13] ), 
        .Y(n2320) );
  AO22X1_LVT U2357 ( .A1(n3364), .A2(wdata[12]), .A3(n3363), .A4(\regs[7][12] ), .Y(n2319) );
  AO22X1_LVT U2358 ( .A1(n3364), .A2(wdata[11]), .A3(n3363), .A4(\regs[7][11] ), .Y(n2318) );
  AO22X1_LVT U2359 ( .A1(n3364), .A2(n3499), .A3(n3363), .A4(\regs[7][10] ), 
        .Y(n2317) );
  AO22X1_LVT U2360 ( .A1(n3364), .A2(wdata[9]), .A3(n3363), .A4(\regs[7][9] ), 
        .Y(n2316) );
  AO22X1_LVT U2362 ( .A1(n3366), .A2(wdata[8]), .A3(n3363), .A4(\regs[7][8] ), 
        .Y(n2315) );
  AO22X1_LVT U2363 ( .A1(n3366), .A2(wdata[7]), .A3(n3363), .A4(\regs[7][7] ), 
        .Y(n2314) );
  AO22X1_LVT U2364 ( .A1(n3366), .A2(wdata[6]), .A3(n3363), .A4(\regs[7][6] ), 
        .Y(n2313) );
  AO22X1_LVT U2365 ( .A1(n3366), .A2(wdata[5]), .A3(n3363), .A4(\regs[7][5] ), 
        .Y(n2312) );
  AO22X1_LVT U2366 ( .A1(n3366), .A2(wdata[4]), .A3(n3363), .A4(\regs[7][4] ), 
        .Y(n2311) );
  AO22X1_LVT U2367 ( .A1(n3366), .A2(wdata[3]), .A3(n3363), .A4(\regs[7][3] ), 
        .Y(n2310) );
  AO22X1_LVT U2368 ( .A1(n3366), .A2(wdata[2]), .A3(n3363), .A4(\regs[7][2] ), 
        .Y(n2309) );
  AO22X1_LVT U2370 ( .A1(n3366), .A2(wdata[1]), .A3(n3363), .A4(\regs[7][1] ), 
        .Y(n2308) );
  AO22X1_LVT U2371 ( .A1(n3366), .A2(wdata[0]), .A3(n3363), .A4(\regs[7][0] ), 
        .Y(n2307) );
  AND4X1_LVT U2372 ( .A1(waddr[3]), .A2(we), .A3(n3002), .A4(n3297), .Y(n3067)
         );
  AND2X1_LVT U2373 ( .A1(n3067), .A2(n3298), .Y(n3030) );
  AO22X1_LVT U2379 ( .A1(n3402), .A2(n3486), .A3(n3401), .A4(\regs[8][31] ), 
        .Y(n2306) );
  AO22X1_LVT U2380 ( .A1(n3402), .A2(wdata[30]), .A3(n3401), .A4(\regs[8][30] ), .Y(n2305) );
  AO22X1_LVT U2381 ( .A1(n3402), .A2(n3453), .A3(n3401), .A4(\regs[8][29] ), 
        .Y(n2304) );
  AO22X1_LVT U2382 ( .A1(n3402), .A2(n3500), .A3(n3401), .A4(\regs[8][28] ), 
        .Y(n2303) );
  AO22X1_LVT U2383 ( .A1(n3402), .A2(wdata[27]), .A3(n3401), .A4(\regs[8][27] ), .Y(n2302) );
  AO22X1_LVT U2384 ( .A1(n3402), .A2(n3503), .A3(n3401), .A4(\regs[8][26] ), 
        .Y(n2301) );
  AO22X1_LVT U2385 ( .A1(n3402), .A2(wdata[25]), .A3(n3401), .A4(\regs[8][25] ), .Y(n2300) );
  AO22X1_LVT U2387 ( .A1(n3398), .A2(n3493), .A3(n3397), .A4(\regs[8][24] ), 
        .Y(n2299) );
  AO22X1_LVT U2388 ( .A1(n3398), .A2(n3497), .A3(n3397), .A4(\regs[8][23] ), 
        .Y(n2298) );
  AO22X1_LVT U2389 ( .A1(n3398), .A2(n3494), .A3(n3397), .A4(\regs[8][22] ), 
        .Y(n2297) );
  AO22X1_LVT U2390 ( .A1(n3398), .A2(wdata[21]), .A3(n3397), .A4(\regs[8][21] ), .Y(n2296) );
  AO22X1_LVT U2391 ( .A1(n3398), .A2(n3469), .A3(n3397), .A4(\regs[8][20] ), 
        .Y(n2295) );
  AO22X1_LVT U2392 ( .A1(n3398), .A2(n3496), .A3(n3397), .A4(\regs[8][19] ), 
        .Y(n2294) );
  AO22X1_LVT U2393 ( .A1(n3398), .A2(n3491), .A3(n3397), .A4(\regs[8][18] ), 
        .Y(n2293) );
  AO22X1_LVT U2394 ( .A1(n3398), .A2(wdata[17]), .A3(n3397), .A4(\regs[8][17] ), .Y(n2292) );
  AO22X1_LVT U2396 ( .A1(n3400), .A2(wdata[16]), .A3(n3399), .A4(\regs[8][16] ), .Y(n2291) );
  AO22X1_LVT U2397 ( .A1(n3400), .A2(n3495), .A3(n3399), .A4(\regs[8][15] ), 
        .Y(n2290) );
  AO22X1_LVT U2398 ( .A1(n3400), .A2(n3498), .A3(n3399), .A4(\regs[8][14] ), 
        .Y(n2289) );
  AO22X1_LVT U2399 ( .A1(n3400), .A2(n3502), .A3(n3399), .A4(\regs[8][13] ), 
        .Y(n2288) );
  AO22X1_LVT U2400 ( .A1(n3402), .A2(wdata[12]), .A3(n3401), .A4(\regs[8][12] ), .Y(n2287) );
  AO22X1_LVT U2401 ( .A1(n3400), .A2(wdata[11]), .A3(n3399), .A4(\regs[8][11] ), .Y(n2286) );
  AO22X1_LVT U2402 ( .A1(n3400), .A2(n3499), .A3(n3399), .A4(\regs[8][10] ), 
        .Y(n2285) );
  AO22X1_LVT U2403 ( .A1(n3402), .A2(wdata[9]), .A3(n3401), .A4(\regs[8][9] ), 
        .Y(n2284) );
  AO22X1_LVT U2405 ( .A1(n3398), .A2(wdata[8]), .A3(n3397), .A4(\regs[8][8] ), 
        .Y(n2283) );
  AO22X1_LVT U2406 ( .A1(n3398), .A2(wdata[7]), .A3(n3397), .A4(\regs[8][7] ), 
        .Y(n2282) );
  AO22X1_LVT U2407 ( .A1(n3398), .A2(wdata[6]), .A3(n3397), .A4(\regs[8][6] ), 
        .Y(n2281) );
  AO22X1_LVT U2408 ( .A1(n3398), .A2(wdata[5]), .A3(n3397), .A4(\regs[8][5] ), 
        .Y(n2280) );
  AO22X1_LVT U2409 ( .A1(n3398), .A2(wdata[4]), .A3(n3397), .A4(\regs[8][4] ), 
        .Y(n2279) );
  AO22X1_LVT U2410 ( .A1(n3398), .A2(wdata[3]), .A3(n3397), .A4(\regs[8][3] ), 
        .Y(n2278) );
  AO22X1_LVT U2411 ( .A1(n3398), .A2(wdata[2]), .A3(n3397), .A4(\regs[8][2] ), 
        .Y(n2277) );
  AO22X1_LVT U2413 ( .A1(n3398), .A2(wdata[1]), .A3(n3397), .A4(\regs[8][1] ), 
        .Y(n2276) );
  AO22X1_LVT U2414 ( .A1(n3398), .A2(wdata[0]), .A3(n3397), .A4(\regs[8][0] ), 
        .Y(n2275) );
  NAND2X0_LVT U2415 ( .A1(n3202), .A2(n3030), .Y(n3012) );
  AO22X1_LVT U2420 ( .A1(n3429), .A2(n3486), .A3(n3428), .A4(\regs[9][31] ), 
        .Y(n2274) );
  AO22X1_LVT U2421 ( .A1(n3429), .A2(wdata[30]), .A3(n3428), .A4(\regs[9][30] ), .Y(n2273) );
  AO22X1_LVT U2422 ( .A1(n3429), .A2(n3501), .A3(n3428), .A4(\regs[9][29] ), 
        .Y(n2272) );
  AO22X1_LVT U2423 ( .A1(n3429), .A2(n3500), .A3(n3428), .A4(\regs[9][28] ), 
        .Y(n2271) );
  AO22X1_LVT U2424 ( .A1(n3429), .A2(wdata[27]), .A3(n3428), .A4(\regs[9][27] ), .Y(n2270) );
  AO22X1_LVT U2425 ( .A1(n3429), .A2(n3503), .A3(n3428), .A4(\regs[9][26] ), 
        .Y(n2269) );
  AO22X1_LVT U2426 ( .A1(n3429), .A2(wdata[25]), .A3(n3428), .A4(\regs[9][25] ), .Y(n2268) );
  AO22X1_LVT U2428 ( .A1(n3431), .A2(n3493), .A3(n3430), .A4(\regs[9][24] ), 
        .Y(n2267) );
  AO22X1_LVT U2429 ( .A1(n3431), .A2(n3497), .A3(n3430), .A4(\regs[9][23] ), 
        .Y(n2266) );
  AO22X1_LVT U2430 ( .A1(n3431), .A2(n3494), .A3(n3430), .A4(\regs[9][22] ), 
        .Y(n2265) );
  AO22X1_LVT U2431 ( .A1(n3431), .A2(wdata[21]), .A3(n3430), .A4(\regs[9][21] ), .Y(n2264) );
  AO22X1_LVT U2432 ( .A1(n3431), .A2(n3483), .A3(n3430), .A4(\regs[9][20] ), 
        .Y(n2263) );
  AO22X1_LVT U2433 ( .A1(n3431), .A2(n3496), .A3(n3430), .A4(\regs[9][19] ), 
        .Y(n2262) );
  AO22X1_LVT U2434 ( .A1(n3431), .A2(n3491), .A3(n3430), .A4(\regs[9][18] ), 
        .Y(n2261) );
  AO22X1_LVT U2435 ( .A1(n3431), .A2(wdata[17]), .A3(n3430), .A4(\regs[9][17] ), .Y(n2260) );
  AO22X1_LVT U2437 ( .A1(n3429), .A2(wdata[16]), .A3(n3428), .A4(\regs[9][16] ), .Y(n2259) );
  AO22X1_LVT U2438 ( .A1(n3429), .A2(n3495), .A3(n3428), .A4(\regs[9][15] ), 
        .Y(n2258) );
  AO22X1_LVT U2439 ( .A1(n3429), .A2(n3498), .A3(n3428), .A4(\regs[9][14] ), 
        .Y(n2257) );
  AO22X1_LVT U2440 ( .A1(n3429), .A2(n3502), .A3(n3428), .A4(\regs[9][13] ), 
        .Y(n2256) );
  AO22X1_LVT U2441 ( .A1(n3429), .A2(wdata[12]), .A3(n3428), .A4(\regs[9][12] ), .Y(n2255) );
  AO22X1_LVT U2442 ( .A1(n3429), .A2(wdata[11]), .A3(n3428), .A4(\regs[9][11] ), .Y(n2254) );
  AO22X1_LVT U2443 ( .A1(n3429), .A2(n3499), .A3(n3428), .A4(\regs[9][10] ), 
        .Y(n2253) );
  AO22X1_LVT U2444 ( .A1(n3429), .A2(wdata[9]), .A3(n3428), .A4(\regs[9][9] ), 
        .Y(n2252) );
  AO22X1_LVT U2446 ( .A1(n3431), .A2(wdata[8]), .A3(n3430), .A4(\regs[9][8] ), 
        .Y(n2251) );
  AO22X1_LVT U2447 ( .A1(n3431), .A2(wdata[7]), .A3(n3430), .A4(\regs[9][7] ), 
        .Y(n2250) );
  AO22X1_LVT U2448 ( .A1(n3431), .A2(wdata[6]), .A3(n3430), .A4(\regs[9][6] ), 
        .Y(n2249) );
  AO22X1_LVT U2449 ( .A1(n3431), .A2(wdata[5]), .A3(n3430), .A4(\regs[9][5] ), 
        .Y(n2248) );
  AO22X1_LVT U2450 ( .A1(n3431), .A2(wdata[4]), .A3(n3430), .A4(\regs[9][4] ), 
        .Y(n2247) );
  AO22X1_LVT U2451 ( .A1(n3431), .A2(wdata[3]), .A3(n3430), .A4(\regs[9][3] ), 
        .Y(n2246) );
  AO22X1_LVT U2452 ( .A1(n3431), .A2(wdata[2]), .A3(n3430), .A4(\regs[9][2] ), 
        .Y(n2245) );
  AO22X1_LVT U2454 ( .A1(n3431), .A2(wdata[1]), .A3(n3430), .A4(\regs[9][1] ), 
        .Y(n2244) );
  AO22X1_LVT U2455 ( .A1(n3431), .A2(wdata[0]), .A3(n3430), .A4(\regs[9][0] ), 
        .Y(n2243) );
  AO22X1_LVT U2461 ( .A1(n3427), .A2(n3486), .A3(n3426), .A4(\regs[10][31] ), 
        .Y(n2242) );
  AO22X1_LVT U2462 ( .A1(n3427), .A2(wdata[30]), .A3(n3426), .A4(
        \regs[10][30] ), .Y(n2241) );
  AO22X1_LVT U2463 ( .A1(n3427), .A2(n3501), .A3(n3426), .A4(\regs[10][29] ), 
        .Y(n2240) );
  AO22X1_LVT U2464 ( .A1(n3427), .A2(n3500), .A3(n3426), .A4(\regs[10][28] ), 
        .Y(n2239) );
  AO22X1_LVT U2465 ( .A1(n3427), .A2(wdata[27]), .A3(n3426), .A4(
        \regs[10][27] ), .Y(n2238) );
  AO22X1_LVT U2466 ( .A1(n3427), .A2(n3503), .A3(n3426), .A4(\regs[10][26] ), 
        .Y(n2237) );
  AO22X1_LVT U2467 ( .A1(n3427), .A2(wdata[25]), .A3(n3426), .A4(
        \regs[10][25] ), .Y(n2236) );
  AO22X1_LVT U2469 ( .A1(n3423), .A2(n3493), .A3(n3021), .A4(\regs[10][24] ), 
        .Y(n2235) );
  AO22X1_LVT U2470 ( .A1(n3425), .A2(n3497), .A3(n3424), .A4(\regs[10][23] ), 
        .Y(n2234) );
  AO22X1_LVT U2471 ( .A1(n3425), .A2(n3494), .A3(n3424), .A4(\regs[10][22] ), 
        .Y(n2233) );
  AO22X1_LVT U2472 ( .A1(n3425), .A2(wdata[21]), .A3(n3424), .A4(
        \regs[10][21] ), .Y(n2232) );
  AO22X1_LVT U2473 ( .A1(n3425), .A2(n3483), .A3(n3424), .A4(\regs[10][20] ), 
        .Y(n2231) );
  AO22X1_LVT U2474 ( .A1(n3425), .A2(n3496), .A3(n3424), .A4(\regs[10][19] ), 
        .Y(n2230) );
  AO22X1_LVT U2475 ( .A1(n3425), .A2(n3491), .A3(n3424), .A4(\regs[10][18] ), 
        .Y(n2229) );
  AO22X1_LVT U2476 ( .A1(n3423), .A2(wdata[17]), .A3(n3021), .A4(
        \regs[10][17] ), .Y(n2228) );
  AO22X1_LVT U2478 ( .A1(n3427), .A2(wdata[16]), .A3(n3426), .A4(
        \regs[10][16] ), .Y(n2227) );
  AO22X1_LVT U2479 ( .A1(n3427), .A2(n3495), .A3(n3426), .A4(\regs[10][15] ), 
        .Y(n2226) );
  AO22X1_LVT U2480 ( .A1(n3427), .A2(n3498), .A3(n3426), .A4(\regs[10][14] ), 
        .Y(n2225) );
  AO22X1_LVT U2481 ( .A1(n3427), .A2(n3502), .A3(n3426), .A4(\regs[10][13] ), 
        .Y(n2224) );
  AO22X1_LVT U2482 ( .A1(n3427), .A2(wdata[12]), .A3(n3426), .A4(
        \regs[10][12] ), .Y(n2223) );
  AO22X1_LVT U2483 ( .A1(n3427), .A2(wdata[11]), .A3(n3426), .A4(
        \regs[10][11] ), .Y(n2222) );
  AO22X1_LVT U2484 ( .A1(n3427), .A2(n3499), .A3(n3426), .A4(\regs[10][10] ), 
        .Y(n2221) );
  AO22X1_LVT U2485 ( .A1(n3427), .A2(wdata[9]), .A3(n3426), .A4(\regs[10][9] ), 
        .Y(n2220) );
  AO22X1_LVT U2487 ( .A1(n3425), .A2(wdata[8]), .A3(n3424), .A4(\regs[10][8] ), 
        .Y(n2219) );
  AO22X1_LVT U2488 ( .A1(n3425), .A2(wdata[7]), .A3(n3424), .A4(\regs[10][7] ), 
        .Y(n2218) );
  AO22X1_LVT U2489 ( .A1(n3425), .A2(wdata[6]), .A3(n3424), .A4(\regs[10][6] ), 
        .Y(n2217) );
  AO22X1_LVT U2490 ( .A1(n3425), .A2(wdata[5]), .A3(n3424), .A4(\regs[10][5] ), 
        .Y(n2216) );
  AO22X1_LVT U2491 ( .A1(n3425), .A2(wdata[4]), .A3(n3424), .A4(\regs[10][4] ), 
        .Y(n2215) );
  AO22X1_LVT U2492 ( .A1(n3425), .A2(wdata[3]), .A3(n3424), .A4(\regs[10][3] ), 
        .Y(n2214) );
  AO22X1_LVT U2493 ( .A1(n3425), .A2(wdata[2]), .A3(n3424), .A4(\regs[10][2] ), 
        .Y(n2213) );
  AO22X1_LVT U2495 ( .A1(n3425), .A2(wdata[1]), .A3(n3424), .A4(\regs[10][1] ), 
        .Y(n2212) );
  AO22X1_LVT U2496 ( .A1(n3425), .A2(wdata[0]), .A3(n3424), .A4(\regs[10][0] ), 
        .Y(n2211) );
  AO22X1_LVT U2502 ( .A1(n3418), .A2(n3486), .A3(n3417), .A4(\regs[11][31] ), 
        .Y(n2210) );
  AO22X1_LVT U2503 ( .A1(n3418), .A2(wdata[30]), .A3(n3417), .A4(
        \regs[11][30] ), .Y(n2209) );
  AO22X1_LVT U2504 ( .A1(n3418), .A2(n3501), .A3(n3417), .A4(\regs[11][29] ), 
        .Y(n2208) );
  AO22X1_LVT U2505 ( .A1(n3418), .A2(n3500), .A3(n3417), .A4(\regs[11][28] ), 
        .Y(n2207) );
  AO22X1_LVT U2506 ( .A1(n3418), .A2(wdata[27]), .A3(n3417), .A4(
        \regs[11][27] ), .Y(n2206) );
  AO22X1_LVT U2507 ( .A1(n3418), .A2(n3503), .A3(n3417), .A4(\regs[11][26] ), 
        .Y(n2205) );
  AO22X1_LVT U2508 ( .A1(n3418), .A2(wdata[25]), .A3(n3417), .A4(
        \regs[11][25] ), .Y(n2204) );
  AO22X1_LVT U2510 ( .A1(n3422), .A2(n3493), .A3(n3421), .A4(\regs[11][24] ), 
        .Y(n2203) );
  AO22X1_LVT U2511 ( .A1(n3420), .A2(n3497), .A3(n3419), .A4(\regs[11][23] ), 
        .Y(n2202) );
  AO22X1_LVT U2512 ( .A1(n3420), .A2(n3494), .A3(n3419), .A4(\regs[11][22] ), 
        .Y(n2201) );
  AO22X1_LVT U2513 ( .A1(n3422), .A2(wdata[21]), .A3(n3421), .A4(
        \regs[11][21] ), .Y(n2200) );
  AO22X1_LVT U2514 ( .A1(n3420), .A2(n3483), .A3(n3419), .A4(\regs[11][20] ), 
        .Y(n2199) );
  AO22X1_LVT U2515 ( .A1(n3422), .A2(n3496), .A3(n3421), .A4(\regs[11][19] ), 
        .Y(n2198) );
  AO22X1_LVT U2516 ( .A1(n3422), .A2(n3491), .A3(n3421), .A4(\regs[11][18] ), 
        .Y(n2197) );
  AO22X1_LVT U2517 ( .A1(n3420), .A2(wdata[17]), .A3(n3419), .A4(
        \regs[11][17] ), .Y(n2196) );
  AO22X1_LVT U2519 ( .A1(n3418), .A2(wdata[16]), .A3(n3417), .A4(
        \regs[11][16] ), .Y(n2195) );
  AO22X1_LVT U2520 ( .A1(n3418), .A2(n3495), .A3(n3417), .A4(\regs[11][15] ), 
        .Y(n2194) );
  AO22X1_LVT U2521 ( .A1(n3418), .A2(n3498), .A3(n3417), .A4(\regs[11][14] ), 
        .Y(n2193) );
  AO22X1_LVT U2522 ( .A1(n3418), .A2(n3502), .A3(n3417), .A4(\regs[11][13] ), 
        .Y(n2192) );
  AO22X1_LVT U2523 ( .A1(n3418), .A2(wdata[12]), .A3(n3417), .A4(
        \regs[11][12] ), .Y(n2191) );
  AO22X1_LVT U2524 ( .A1(n3418), .A2(wdata[11]), .A3(n3417), .A4(
        \regs[11][11] ), .Y(n2190) );
  AO22X1_LVT U2525 ( .A1(n3418), .A2(n3499), .A3(n3417), .A4(\regs[11][10] ), 
        .Y(n2189) );
  AO22X1_LVT U2526 ( .A1(n3418), .A2(wdata[9]), .A3(n3417), .A4(\regs[11][9] ), 
        .Y(n2188) );
  AO22X1_LVT U2528 ( .A1(n3422), .A2(wdata[8]), .A3(n3421), .A4(\regs[11][8] ), 
        .Y(n2187) );
  AO22X1_LVT U2529 ( .A1(n3420), .A2(wdata[7]), .A3(n3419), .A4(\regs[11][7] ), 
        .Y(n2186) );
  AO22X1_LVT U2530 ( .A1(n3420), .A2(wdata[6]), .A3(n3419), .A4(\regs[11][6] ), 
        .Y(n2185) );
  AO22X1_LVT U2531 ( .A1(n3420), .A2(wdata[5]), .A3(n3419), .A4(\regs[11][5] ), 
        .Y(n2184) );
  AO22X1_LVT U2532 ( .A1(n3422), .A2(wdata[4]), .A3(n3421), .A4(\regs[11][4] ), 
        .Y(n2183) );
  AO22X1_LVT U2533 ( .A1(n3422), .A2(wdata[3]), .A3(n3421), .A4(\regs[11][3] ), 
        .Y(n2182) );
  AO22X1_LVT U2534 ( .A1(n3420), .A2(wdata[2]), .A3(n3419), .A4(\regs[11][2] ), 
        .Y(n2181) );
  AO22X1_LVT U2536 ( .A1(n3420), .A2(wdata[1]), .A3(n3419), .A4(\regs[11][1] ), 
        .Y(n2180) );
  AO22X1_LVT U2537 ( .A1(n3420), .A2(wdata[0]), .A3(n3419), .A4(\regs[11][0] ), 
        .Y(n2179) );
  NAND4X0_LVT U2538 ( .A1(n3470), .A2(n3067), .A3(n3192), .A4(n3191), .Y(n3040) );
  AO22X1_LVT U2543 ( .A1(n3312), .A2(n3486), .A3(n3311), .A4(\regs[12][31] ), 
        .Y(n2178) );
  AO22X1_LVT U2544 ( .A1(n3312), .A2(wdata[30]), .A3(n3311), .A4(
        \regs[12][30] ), .Y(n2177) );
  AO22X1_LVT U2545 ( .A1(n3312), .A2(n3501), .A3(n3311), .A4(\regs[12][29] ), 
        .Y(n2176) );
  AO22X1_LVT U2546 ( .A1(n3312), .A2(n3500), .A3(n3311), .A4(\regs[12][28] ), 
        .Y(n2175) );
  AO22X1_LVT U2547 ( .A1(n3312), .A2(wdata[27]), .A3(n3311), .A4(
        \regs[12][27] ), .Y(n2174) );
  AO22X1_LVT U2548 ( .A1(n3312), .A2(n3503), .A3(n3311), .A4(\regs[12][26] ), 
        .Y(n2173) );
  AO22X1_LVT U2549 ( .A1(n3312), .A2(wdata[25]), .A3(n3311), .A4(
        \regs[12][25] ), .Y(n2172) );
  AO22X1_LVT U2551 ( .A1(n3314), .A2(n3493), .A3(n3313), .A4(\regs[12][24] ), 
        .Y(n2171) );
  AO22X1_LVT U2552 ( .A1(n3312), .A2(n3497), .A3(n3311), .A4(\regs[12][23] ), 
        .Y(n2170) );
  AO22X1_LVT U2553 ( .A1(n3312), .A2(n3494), .A3(n3311), .A4(\regs[12][22] ), 
        .Y(n2169) );
  AO22X1_LVT U2554 ( .A1(n3314), .A2(wdata[21]), .A3(n3313), .A4(
        \regs[12][21] ), .Y(n2168) );
  AO22X1_LVT U2555 ( .A1(n3312), .A2(n3483), .A3(n3311), .A4(\regs[12][20] ), 
        .Y(n2167) );
  AO22X1_LVT U2556 ( .A1(n3312), .A2(n3496), .A3(n3311), .A4(\regs[12][19] ), 
        .Y(n2166) );
  AO22X1_LVT U2557 ( .A1(n3312), .A2(n3491), .A3(n3311), .A4(\regs[12][18] ), 
        .Y(n2165) );
  AO22X1_LVT U2558 ( .A1(n3314), .A2(wdata[17]), .A3(n3313), .A4(
        \regs[12][17] ), .Y(n2164) );
  AO22X1_LVT U2560 ( .A1(n3312), .A2(wdata[16]), .A3(n3311), .A4(
        \regs[12][16] ), .Y(n2163) );
  AO22X1_LVT U2561 ( .A1(n3312), .A2(n3495), .A3(n3311), .A4(\regs[12][15] ), 
        .Y(n2162) );
  AO22X1_LVT U2562 ( .A1(n3312), .A2(n3498), .A3(n3311), .A4(\regs[12][14] ), 
        .Y(n2161) );
  AO22X1_LVT U2563 ( .A1(n3312), .A2(n3502), .A3(n3311), .A4(\regs[12][13] ), 
        .Y(n2160) );
  AO22X1_LVT U2564 ( .A1(n3312), .A2(wdata[12]), .A3(n3311), .A4(
        \regs[12][12] ), .Y(n2159) );
  AO22X1_LVT U2565 ( .A1(n3312), .A2(wdata[11]), .A3(n3311), .A4(
        \regs[12][11] ), .Y(n2158) );
  AO22X1_LVT U2566 ( .A1(n3312), .A2(n3499), .A3(n3311), .A4(\regs[12][10] ), 
        .Y(n2157) );
  AO22X1_LVT U2567 ( .A1(n3312), .A2(wdata[9]), .A3(n3311), .A4(\regs[12][9] ), 
        .Y(n2156) );
  AO22X1_LVT U2569 ( .A1(n3314), .A2(wdata[8]), .A3(n3313), .A4(\regs[12][8] ), 
        .Y(n2155) );
  AO22X1_LVT U2570 ( .A1(n3314), .A2(wdata[7]), .A3(n3313), .A4(\regs[12][7] ), 
        .Y(n2154) );
  AO22X1_LVT U2571 ( .A1(n3314), .A2(wdata[6]), .A3(n3313), .A4(\regs[12][6] ), 
        .Y(n2153) );
  AO22X1_LVT U2572 ( .A1(n3314), .A2(wdata[5]), .A3(n3313), .A4(\regs[12][5] ), 
        .Y(n2152) );
  AO22X1_LVT U2573 ( .A1(n3314), .A2(wdata[4]), .A3(n3313), .A4(\regs[12][4] ), 
        .Y(n2151) );
  AO22X1_LVT U2574 ( .A1(n3314), .A2(wdata[3]), .A3(n3313), .A4(\regs[12][3] ), 
        .Y(n2150) );
  AO22X1_LVT U2575 ( .A1(n3314), .A2(wdata[2]), .A3(n3313), .A4(\regs[12][2] ), 
        .Y(n2149) );
  AO22X1_LVT U2577 ( .A1(n3314), .A2(wdata[1]), .A3(n3313), .A4(\regs[12][1] ), 
        .Y(n2148) );
  AO22X1_LVT U2578 ( .A1(n3314), .A2(wdata[0]), .A3(n3313), .A4(\regs[12][0] ), 
        .Y(n2147) );
  NAND3X0_LVT U2579 ( .A1(n3470), .A2(n3202), .A3(n3067), .Y(n3049) );
  AO22X1_LVT U2584 ( .A1(n3359), .A2(n3486), .A3(n3358), .A4(\regs[13][31] ), 
        .Y(n2146) );
  AO22X1_LVT U2585 ( .A1(n3359), .A2(wdata[30]), .A3(n3358), .A4(
        \regs[13][30] ), .Y(n2145) );
  AO22X1_LVT U2586 ( .A1(n3359), .A2(n3501), .A3(n3358), .A4(\regs[13][29] ), 
        .Y(n2144) );
  AO22X1_LVT U2587 ( .A1(n3359), .A2(n3500), .A3(n3358), .A4(\regs[13][28] ), 
        .Y(n2143) );
  AO22X1_LVT U2588 ( .A1(n3359), .A2(wdata[27]), .A3(n3358), .A4(
        \regs[13][27] ), .Y(n2142) );
  AO22X1_LVT U2589 ( .A1(n3359), .A2(n3503), .A3(n3358), .A4(\regs[13][26] ), 
        .Y(n2141) );
  AO22X1_LVT U2590 ( .A1(n3359), .A2(wdata[25]), .A3(n3358), .A4(
        \regs[13][25] ), .Y(n2140) );
  AO22X1_LVT U2592 ( .A1(n3359), .A2(n3493), .A3(n3358), .A4(\regs[13][24] ), 
        .Y(n2139) );
  AO22X1_LVT U2593 ( .A1(n3359), .A2(n3497), .A3(n3358), .A4(\regs[13][23] ), 
        .Y(n2138) );
  AO22X1_LVT U2594 ( .A1(n3361), .A2(n3494), .A3(n3360), .A4(\regs[13][22] ), 
        .Y(n2137) );
  AO22X1_LVT U2595 ( .A1(n3359), .A2(wdata[21]), .A3(n3358), .A4(
        \regs[13][21] ), .Y(n2136) );
  AO22X1_LVT U2596 ( .A1(n3361), .A2(n3483), .A3(n3360), .A4(\regs[13][20] ), 
        .Y(n2135) );
  AO22X1_LVT U2597 ( .A1(n3361), .A2(n3496), .A3(n3360), .A4(\regs[13][19] ), 
        .Y(n2134) );
  AO22X1_LVT U2598 ( .A1(n3361), .A2(n3491), .A3(n3360), .A4(\regs[13][18] ), 
        .Y(n2133) );
  AO22X1_LVT U2599 ( .A1(n3359), .A2(wdata[17]), .A3(n3358), .A4(
        \regs[13][17] ), .Y(n2132) );
  AO22X1_LVT U2601 ( .A1(n3359), .A2(wdata[16]), .A3(n3358), .A4(
        \regs[13][16] ), .Y(n2131) );
  AO22X1_LVT U2602 ( .A1(n3359), .A2(n3495), .A3(n3358), .A4(\regs[13][15] ), 
        .Y(n2130) );
  AO22X1_LVT U2603 ( .A1(n3359), .A2(n3498), .A3(n3358), .A4(\regs[13][14] ), 
        .Y(n2129) );
  AO22X1_LVT U2604 ( .A1(n3359), .A2(n3502), .A3(n3358), .A4(\regs[13][13] ), 
        .Y(n2128) );
  AO22X1_LVT U2605 ( .A1(n3359), .A2(wdata[12]), .A3(n3358), .A4(
        \regs[13][12] ), .Y(n2127) );
  AO22X1_LVT U2606 ( .A1(n3359), .A2(wdata[11]), .A3(n3358), .A4(
        \regs[13][11] ), .Y(n2126) );
  AO22X1_LVT U2607 ( .A1(n3359), .A2(wdata[10]), .A3(n3358), .A4(
        \regs[13][10] ), .Y(n2125) );
  AO22X1_LVT U2608 ( .A1(n3359), .A2(wdata[9]), .A3(n3358), .A4(\regs[13][9] ), 
        .Y(n2124) );
  AO22X1_LVT U2610 ( .A1(n3361), .A2(wdata[8]), .A3(n3360), .A4(\regs[13][8] ), 
        .Y(n2123) );
  AO22X1_LVT U2611 ( .A1(n3361), .A2(wdata[7]), .A3(n3360), .A4(\regs[13][7] ), 
        .Y(n2122) );
  AO22X1_LVT U2612 ( .A1(n3361), .A2(wdata[6]), .A3(n3360), .A4(\regs[13][6] ), 
        .Y(n2121) );
  AO22X1_LVT U2613 ( .A1(n3361), .A2(wdata[5]), .A3(n3360), .A4(\regs[13][5] ), 
        .Y(n2120) );
  AO22X1_LVT U2614 ( .A1(n3361), .A2(wdata[4]), .A3(n3360), .A4(\regs[13][4] ), 
        .Y(n2119) );
  AO22X1_LVT U2615 ( .A1(n3361), .A2(wdata[3]), .A3(n3360), .A4(\regs[13][3] ), 
        .Y(n2118) );
  AO22X1_LVT U2616 ( .A1(n3361), .A2(wdata[2]), .A3(n3360), .A4(\regs[13][2] ), 
        .Y(n2117) );
  AO22X1_LVT U2618 ( .A1(n3361), .A2(wdata[1]), .A3(n3360), .A4(\regs[13][1] ), 
        .Y(n2116) );
  AO22X1_LVT U2619 ( .A1(n3361), .A2(wdata[0]), .A3(n3360), .A4(\regs[13][0] ), 
        .Y(n2115) );
  AO22X1_LVT U2625 ( .A1(n3353), .A2(n3486), .A3(n3352), .A4(\regs[14][31] ), 
        .Y(n2114) );
  AO22X1_LVT U2626 ( .A1(n3353), .A2(wdata[30]), .A3(n3352), .A4(
        \regs[14][30] ), .Y(n2113) );
  AO22X1_LVT U2627 ( .A1(n3353), .A2(n3501), .A3(n3352), .A4(\regs[14][29] ), 
        .Y(n2112) );
  AO22X1_LVT U2628 ( .A1(n3353), .A2(n3500), .A3(n3352), .A4(\regs[14][28] ), 
        .Y(n2111) );
  AO22X1_LVT U2629 ( .A1(n3353), .A2(wdata[27]), .A3(n3352), .A4(
        \regs[14][27] ), .Y(n2110) );
  AO22X1_LVT U2630 ( .A1(n3353), .A2(n3503), .A3(n3352), .A4(\regs[14][26] ), 
        .Y(n2109) );
  AO22X1_LVT U2631 ( .A1(n3353), .A2(wdata[25]), .A3(n3352), .A4(
        \regs[14][25] ), .Y(n2108) );
  AO22X1_LVT U2633 ( .A1(n3353), .A2(n3493), .A3(n3352), .A4(\regs[14][24] ), 
        .Y(n2107) );
  AO22X1_LVT U2634 ( .A1(n3353), .A2(n3497), .A3(n3352), .A4(\regs[14][23] ), 
        .Y(n2106) );
  AO22X1_LVT U2635 ( .A1(n3353), .A2(n3494), .A3(n3352), .A4(\regs[14][22] ), 
        .Y(n2105) );
  AO22X1_LVT U2636 ( .A1(n3353), .A2(wdata[21]), .A3(n3352), .A4(
        \regs[14][21] ), .Y(n2104) );
  AO22X1_LVT U2637 ( .A1(n3353), .A2(n3483), .A3(n3352), .A4(\regs[14][20] ), 
        .Y(n2103) );
  AO22X1_LVT U2638 ( .A1(n3353), .A2(n3496), .A3(n3352), .A4(\regs[14][19] ), 
        .Y(n2102) );
  AO22X1_LVT U2639 ( .A1(n3353), .A2(n3491), .A3(n3352), .A4(\regs[14][18] ), 
        .Y(n2101) );
  AO22X1_LVT U2640 ( .A1(n3357), .A2(wdata[17]), .A3(n3356), .A4(
        \regs[14][17] ), .Y(n2100) );
  AO22X1_LVT U2642 ( .A1(n3355), .A2(wdata[16]), .A3(n3354), .A4(
        \regs[14][16] ), .Y(n2099) );
  AO22X1_LVT U2643 ( .A1(n3355), .A2(n3495), .A3(n3354), .A4(\regs[14][15] ), 
        .Y(n2098) );
  AO22X1_LVT U2644 ( .A1(n3353), .A2(n3498), .A3(n3352), .A4(\regs[14][14] ), 
        .Y(n2097) );
  AO22X1_LVT U2645 ( .A1(n3355), .A2(n3502), .A3(n3354), .A4(\regs[14][13] ), 
        .Y(n2096) );
  AO22X1_LVT U2646 ( .A1(n3355), .A2(wdata[12]), .A3(n3354), .A4(
        \regs[14][12] ), .Y(n2095) );
  AO22X1_LVT U2647 ( .A1(n3353), .A2(wdata[11]), .A3(n3352), .A4(
        \regs[14][11] ), .Y(n2094) );
  AO22X1_LVT U2648 ( .A1(n3355), .A2(n3499), .A3(n3354), .A4(\regs[14][10] ), 
        .Y(n2093) );
  AO22X1_LVT U2649 ( .A1(n3355), .A2(wdata[9]), .A3(n3354), .A4(\regs[14][9] ), 
        .Y(n2092) );
  AO22X1_LVT U2651 ( .A1(n3357), .A2(wdata[8]), .A3(n3356), .A4(\regs[14][8] ), 
        .Y(n2091) );
  AO22X1_LVT U2652 ( .A1(n3357), .A2(wdata[7]), .A3(n3356), .A4(\regs[14][7] ), 
        .Y(n2090) );
  AO22X1_LVT U2653 ( .A1(n3357), .A2(wdata[6]), .A3(n3356), .A4(\regs[14][6] ), 
        .Y(n2089) );
  AO22X1_LVT U2654 ( .A1(n3357), .A2(wdata[5]), .A3(n3356), .A4(\regs[14][5] ), 
        .Y(n2088) );
  AO22X1_LVT U2655 ( .A1(n3357), .A2(wdata[4]), .A3(n3356), .A4(\regs[14][4] ), 
        .Y(n2087) );
  AO22X1_LVT U2656 ( .A1(n3357), .A2(wdata[3]), .A3(n3356), .A4(\regs[14][3] ), 
        .Y(n2086) );
  AO22X1_LVT U2657 ( .A1(n3357), .A2(wdata[2]), .A3(n3356), .A4(\regs[14][2] ), 
        .Y(n2085) );
  AO22X1_LVT U2659 ( .A1(n3357), .A2(wdata[1]), .A3(n3356), .A4(\regs[14][1] ), 
        .Y(n2084) );
  AO22X1_LVT U2660 ( .A1(n3357), .A2(wdata[0]), .A3(n3356), .A4(\regs[14][0] ), 
        .Y(n2083) );
  AO22X1_LVT U2666 ( .A1(n3349), .A2(wdata[31]), .A3(n3348), .A4(
        \regs[15][31] ), .Y(n2082) );
  AO22X1_LVT U2667 ( .A1(n3349), .A2(wdata[30]), .A3(n3348), .A4(
        \regs[15][30] ), .Y(n2081) );
  AO22X1_LVT U2668 ( .A1(n3349), .A2(n3501), .A3(n3348), .A4(\regs[15][29] ), 
        .Y(n2080) );
  AO22X1_LVT U2669 ( .A1(n3349), .A2(n3500), .A3(n3348), .A4(\regs[15][28] ), 
        .Y(n2079) );
  AO22X1_LVT U2670 ( .A1(n3349), .A2(wdata[27]), .A3(n3348), .A4(
        \regs[15][27] ), .Y(n2078) );
  AO22X1_LVT U2671 ( .A1(n3349), .A2(n3503), .A3(n3348), .A4(\regs[15][26] ), 
        .Y(n2077) );
  AO22X1_LVT U2672 ( .A1(n3349), .A2(wdata[25]), .A3(n3348), .A4(
        \regs[15][25] ), .Y(n2076) );
  AO22X1_LVT U2674 ( .A1(n3349), .A2(wdata[24]), .A3(n3348), .A4(
        \regs[15][24] ), .Y(n2075) );
  AO22X1_LVT U2675 ( .A1(n3349), .A2(wdata[23]), .A3(n3348), .A4(
        \regs[15][23] ), .Y(n2074) );
  AO22X1_LVT U2676 ( .A1(n3347), .A2(wdata[22]), .A3(n3348), .A4(
        \regs[15][22] ), .Y(n2073) );
  AO22X1_LVT U2677 ( .A1(n3351), .A2(wdata[21]), .A3(n3348), .A4(
        \regs[15][21] ), .Y(n2072) );
  AO22X1_LVT U2678 ( .A1(n3349), .A2(n3492), .A3(n3348), .A4(\regs[15][20] ), 
        .Y(n2071) );
  AO22X1_LVT U2679 ( .A1(n3349), .A2(n3496), .A3(n3348), .A4(\regs[15][19] ), 
        .Y(n2070) );
  AO22X1_LVT U2680 ( .A1(n3347), .A2(wdata[18]), .A3(n3348), .A4(
        \regs[15][18] ), .Y(n2069) );
  AO22X1_LVT U2681 ( .A1(n3351), .A2(wdata[17]), .A3(n3348), .A4(
        \regs[15][17] ), .Y(n2068) );
  AO22X1_LVT U2683 ( .A1(n3349), .A2(wdata[16]), .A3(n3348), .A4(
        \regs[15][16] ), .Y(n2067) );
  AO22X1_LVT U2684 ( .A1(n3349), .A2(wdata[15]), .A3(n3348), .A4(
        \regs[15][15] ), .Y(n2066) );
  AO22X1_LVT U2685 ( .A1(n3349), .A2(n3498), .A3(n3348), .A4(\regs[15][14] ), 
        .Y(n2065) );
  AO22X1_LVT U2686 ( .A1(n3349), .A2(wdata[13]), .A3(n3348), .A4(
        \regs[15][13] ), .Y(n2064) );
  AO22X1_LVT U2687 ( .A1(n3349), .A2(wdata[12]), .A3(n3348), .A4(
        \regs[15][12] ), .Y(n2063) );
  AO22X1_LVT U2688 ( .A1(n3349), .A2(wdata[11]), .A3(n3348), .A4(
        \regs[15][11] ), .Y(n2062) );
  AO22X1_LVT U2689 ( .A1(n3349), .A2(n3499), .A3(n3348), .A4(\regs[15][10] ), 
        .Y(n2061) );
  AO22X1_LVT U2690 ( .A1(n3349), .A2(wdata[9]), .A3(n3348), .A4(\regs[15][9] ), 
        .Y(n2060) );
  AO22X1_LVT U2692 ( .A1(n3351), .A2(wdata[8]), .A3(n3348), .A4(\regs[15][8] ), 
        .Y(n2059) );
  AO22X1_LVT U2693 ( .A1(n3351), .A2(wdata[7]), .A3(n3348), .A4(\regs[15][7] ), 
        .Y(n2058) );
  AO22X1_LVT U2694 ( .A1(n3351), .A2(wdata[6]), .A3(n3348), .A4(\regs[15][6] ), 
        .Y(n2057) );
  AO22X1_LVT U2695 ( .A1(n3351), .A2(wdata[5]), .A3(n3348), .A4(\regs[15][5] ), 
        .Y(n2056) );
  AO22X1_LVT U2696 ( .A1(n3351), .A2(wdata[4]), .A3(n3348), .A4(\regs[15][4] ), 
        .Y(n2055) );
  AO22X1_LVT U2697 ( .A1(n3351), .A2(wdata[3]), .A3(n3348), .A4(\regs[15][3] ), 
        .Y(n2054) );
  AO22X1_LVT U2698 ( .A1(n3351), .A2(wdata[2]), .A3(n3348), .A4(\regs[15][2] ), 
        .Y(n2053) );
  AO22X1_LVT U2700 ( .A1(n3351), .A2(wdata[1]), .A3(n3348), .A4(\regs[15][1] ), 
        .Y(n2052) );
  AO22X1_LVT U2701 ( .A1(n3351), .A2(wdata[0]), .A3(n3348), .A4(\regs[15][0] ), 
        .Y(n2051) );
  AND4X1_LVT U2702 ( .A1(waddr[4]), .A2(we), .A3(n3077), .A4(n3297), .Y(n3142)
         );
  AND2X1_LVT U2703 ( .A1(n3142), .A2(n3298), .Y(n3105) );
  NAND3X0_LVT U2704 ( .A1(n3105), .A2(n3192), .A3(n3191), .Y(n3078) );
  AO22X1_LVT U2709 ( .A1(n3394), .A2(n3486), .A3(n3393), .A4(\regs[16][31] ), 
        .Y(n2050) );
  AO22X1_LVT U2710 ( .A1(n3394), .A2(wdata[30]), .A3(n3393), .A4(
        \regs[16][30] ), .Y(n2049) );
  AO22X1_LVT U2711 ( .A1(n3394), .A2(n3501), .A3(n3393), .A4(\regs[16][29] ), 
        .Y(n2048) );
  AO22X1_LVT U2712 ( .A1(n3394), .A2(n3500), .A3(n3393), .A4(\regs[16][28] ), 
        .Y(n2047) );
  AO22X1_LVT U2713 ( .A1(n3394), .A2(wdata[27]), .A3(n3393), .A4(
        \regs[16][27] ), .Y(n2046) );
  AO22X1_LVT U2714 ( .A1(n3394), .A2(n3503), .A3(n3393), .A4(\regs[16][26] ), 
        .Y(n2045) );
  AO22X1_LVT U2715 ( .A1(n3394), .A2(wdata[25]), .A3(n3393), .A4(
        \regs[16][25] ), .Y(n2044) );
  AO22X1_LVT U2717 ( .A1(n3394), .A2(n3493), .A3(n3393), .A4(\regs[16][24] ), 
        .Y(n2043) );
  AO22X1_LVT U2718 ( .A1(n3394), .A2(n3497), .A3(n3393), .A4(\regs[16][23] ), 
        .Y(n2042) );
  AO22X1_LVT U2719 ( .A1(n3394), .A2(n3494), .A3(n3393), .A4(\regs[16][22] ), 
        .Y(n2041) );
  AO22X1_LVT U2720 ( .A1(n3396), .A2(wdata[21]), .A3(n3395), .A4(
        \regs[16][21] ), .Y(n2040) );
  AO22X1_LVT U2721 ( .A1(n3394), .A2(n3483), .A3(n3393), .A4(\regs[16][20] ), 
        .Y(n2039) );
  AO22X1_LVT U2722 ( .A1(n3396), .A2(n3496), .A3(n3395), .A4(\regs[16][19] ), 
        .Y(n2038) );
  AO22X1_LVT U2723 ( .A1(n3396), .A2(n3491), .A3(n3395), .A4(\regs[16][18] ), 
        .Y(n2037) );
  AO22X1_LVT U2724 ( .A1(n3394), .A2(wdata[17]), .A3(n3393), .A4(
        \regs[16][17] ), .Y(n2036) );
  AO22X1_LVT U2726 ( .A1(n3394), .A2(wdata[16]), .A3(n3393), .A4(
        \regs[16][16] ), .Y(n2035) );
  AO22X1_LVT U2727 ( .A1(n3394), .A2(n3495), .A3(n3393), .A4(\regs[16][15] ), 
        .Y(n2034) );
  AO22X1_LVT U2728 ( .A1(n3394), .A2(n3498), .A3(n3393), .A4(\regs[16][14] ), 
        .Y(n2033) );
  AO22X1_LVT U2729 ( .A1(n3394), .A2(n3502), .A3(n3393), .A4(\regs[16][13] ), 
        .Y(n2032) );
  AO22X1_LVT U2730 ( .A1(n3394), .A2(wdata[12]), .A3(n3393), .A4(
        \regs[16][12] ), .Y(n2031) );
  AO22X1_LVT U2731 ( .A1(n3394), .A2(wdata[11]), .A3(n3393), .A4(
        \regs[16][11] ), .Y(n2030) );
  AO22X1_LVT U2732 ( .A1(n3394), .A2(n3499), .A3(n3393), .A4(\regs[16][10] ), 
        .Y(n2029) );
  AO22X1_LVT U2733 ( .A1(n3394), .A2(wdata[9]), .A3(n3393), .A4(\regs[16][9] ), 
        .Y(n2028) );
  AO22X1_LVT U2735 ( .A1(n3396), .A2(wdata[8]), .A3(n3395), .A4(\regs[16][8] ), 
        .Y(n2027) );
  AO22X1_LVT U2736 ( .A1(n3396), .A2(wdata[7]), .A3(n3395), .A4(\regs[16][7] ), 
        .Y(n2026) );
  AO22X1_LVT U2737 ( .A1(n3396), .A2(wdata[6]), .A3(n3395), .A4(\regs[16][6] ), 
        .Y(n2025) );
  AO22X1_LVT U2738 ( .A1(n3396), .A2(wdata[5]), .A3(n3395), .A4(\regs[16][5] ), 
        .Y(n2024) );
  AO22X1_LVT U2739 ( .A1(n3396), .A2(wdata[4]), .A3(n3395), .A4(\regs[16][4] ), 
        .Y(n2023) );
  AO22X1_LVT U2740 ( .A1(n3396), .A2(wdata[3]), .A3(n3395), .A4(\regs[16][3] ), 
        .Y(n2022) );
  AO22X1_LVT U2741 ( .A1(n3396), .A2(wdata[2]), .A3(n3395), .A4(\regs[16][2] ), 
        .Y(n2021) );
  AO22X1_LVT U2743 ( .A1(n3396), .A2(wdata[1]), .A3(n3395), .A4(\regs[16][1] ), 
        .Y(n2020) );
  AO22X1_LVT U2744 ( .A1(n3396), .A2(wdata[0]), .A3(n3395), .A4(\regs[16][0] ), 
        .Y(n2019) );
  NAND2X0_LVT U2745 ( .A1(n3202), .A2(n3105), .Y(n3087) );
  AO22X1_LVT U2750 ( .A1(n3414), .A2(n3486), .A3(n3413), .A4(\regs[17][31] ), 
        .Y(n2018) );
  AO22X1_LVT U2751 ( .A1(n3414), .A2(wdata[30]), .A3(n3413), .A4(
        \regs[17][30] ), .Y(n2017) );
  AO22X1_LVT U2752 ( .A1(n3414), .A2(n3501), .A3(n3413), .A4(\regs[17][29] ), 
        .Y(n2016) );
  AO22X1_LVT U2753 ( .A1(n3414), .A2(n3500), .A3(n3413), .A4(\regs[17][28] ), 
        .Y(n2015) );
  AO22X1_LVT U2754 ( .A1(n3414), .A2(wdata[27]), .A3(n3413), .A4(
        \regs[17][27] ), .Y(n2014) );
  AO22X1_LVT U2755 ( .A1(n3414), .A2(n3503), .A3(n3413), .A4(\regs[17][26] ), 
        .Y(n2013) );
  AO22X1_LVT U2756 ( .A1(n3414), .A2(wdata[25]), .A3(n3413), .A4(
        \regs[17][25] ), .Y(n2012) );
  AO22X1_LVT U2758 ( .A1(n3416), .A2(n3493), .A3(n3415), .A4(\regs[17][24] ), 
        .Y(n2011) );
  AO22X1_LVT U2759 ( .A1(n3414), .A2(n3497), .A3(n3413), .A4(\regs[17][23] ), 
        .Y(n2010) );
  AO22X1_LVT U2760 ( .A1(n3416), .A2(n3494), .A3(n3415), .A4(\regs[17][22] ), 
        .Y(n2009) );
  AO22X1_LVT U2761 ( .A1(n3416), .A2(wdata[21]), .A3(n3415), .A4(
        \regs[17][21] ), .Y(n2008) );
  AO22X1_LVT U2762 ( .A1(n3414), .A2(n3483), .A3(n3413), .A4(\regs[17][20] ), 
        .Y(n2007) );
  AO22X1_LVT U2763 ( .A1(n3414), .A2(n3496), .A3(n3413), .A4(\regs[17][19] ), 
        .Y(n2006) );
  AO22X1_LVT U2764 ( .A1(n3414), .A2(n3491), .A3(n3413), .A4(\regs[17][18] ), 
        .Y(n2005) );
  AO22X1_LVT U2765 ( .A1(n3416), .A2(wdata[17]), .A3(n3415), .A4(
        \regs[17][17] ), .Y(n2004) );
  AO22X1_LVT U2767 ( .A1(n3414), .A2(wdata[16]), .A3(n3413), .A4(
        \regs[17][16] ), .Y(n2003) );
  AO22X1_LVT U2768 ( .A1(n3414), .A2(n3495), .A3(n3413), .A4(\regs[17][15] ), 
        .Y(n2002) );
  AO22X1_LVT U2769 ( .A1(n3414), .A2(n3498), .A3(n3413), .A4(\regs[17][14] ), 
        .Y(n2001) );
  AO22X1_LVT U2770 ( .A1(n3414), .A2(n3502), .A3(n3413), .A4(\regs[17][13] ), 
        .Y(n2000) );
  AO22X1_LVT U2771 ( .A1(n3414), .A2(wdata[12]), .A3(n3413), .A4(
        \regs[17][12] ), .Y(n1999) );
  AO22X1_LVT U2772 ( .A1(n3414), .A2(wdata[11]), .A3(n3413), .A4(
        \regs[17][11] ), .Y(n1998) );
  AO22X1_LVT U2773 ( .A1(n3414), .A2(n3499), .A3(n3413), .A4(\regs[17][10] ), 
        .Y(n1997) );
  AO22X1_LVT U2774 ( .A1(n3414), .A2(wdata[9]), .A3(n3413), .A4(\regs[17][9] ), 
        .Y(n1996) );
  AO22X1_LVT U2776 ( .A1(n3416), .A2(wdata[8]), .A3(n3415), .A4(\regs[17][8] ), 
        .Y(n1995) );
  AO22X1_LVT U2777 ( .A1(n3416), .A2(wdata[7]), .A3(n3415), .A4(\regs[17][7] ), 
        .Y(n1994) );
  AO22X1_LVT U2778 ( .A1(n3416), .A2(wdata[6]), .A3(n3415), .A4(\regs[17][6] ), 
        .Y(n1993) );
  AO22X1_LVT U2779 ( .A1(n3416), .A2(wdata[5]), .A3(n3415), .A4(\regs[17][5] ), 
        .Y(n1992) );
  AO22X1_LVT U2780 ( .A1(n3416), .A2(wdata[4]), .A3(n3415), .A4(\regs[17][4] ), 
        .Y(n1991) );
  AO22X1_LVT U2781 ( .A1(n3416), .A2(wdata[3]), .A3(n3415), .A4(\regs[17][3] ), 
        .Y(n1990) );
  AO22X1_LVT U2782 ( .A1(n3416), .A2(wdata[2]), .A3(n3415), .A4(\regs[17][2] ), 
        .Y(n1989) );
  AO22X1_LVT U2784 ( .A1(n3416), .A2(wdata[1]), .A3(n3415), .A4(\regs[17][1] ), 
        .Y(n1988) );
  AO22X1_LVT U2785 ( .A1(n3416), .A2(wdata[0]), .A3(n3415), .A4(\regs[17][0] ), 
        .Y(n1987) );
  AO22X1_LVT U2791 ( .A1(n3410), .A2(n3486), .A3(n3409), .A4(\regs[18][31] ), 
        .Y(n1986) );
  AO22X1_LVT U2792 ( .A1(n3410), .A2(wdata[30]), .A3(n3409), .A4(
        \regs[18][30] ), .Y(n1985) );
  AO22X1_LVT U2793 ( .A1(n3412), .A2(n3501), .A3(n3411), .A4(\regs[18][29] ), 
        .Y(n1984) );
  AO22X1_LVT U2794 ( .A1(n3412), .A2(n3500), .A3(n3411), .A4(\regs[18][28] ), 
        .Y(n1983) );
  AO22X1_LVT U2795 ( .A1(n3412), .A2(wdata[27]), .A3(n3411), .A4(
        \regs[18][27] ), .Y(n1982) );
  AO22X1_LVT U2796 ( .A1(n3412), .A2(n3503), .A3(n3411), .A4(\regs[18][26] ), 
        .Y(n1981) );
  AO22X1_LVT U2797 ( .A1(n3410), .A2(wdata[25]), .A3(n3409), .A4(
        \regs[18][25] ), .Y(n1980) );
  AO22X1_LVT U2799 ( .A1(n3410), .A2(n3493), .A3(n3409), .A4(\regs[18][24] ), 
        .Y(n1979) );
  AO22X1_LVT U2800 ( .A1(n3412), .A2(n3497), .A3(n3411), .A4(\regs[18][23] ), 
        .Y(n1978) );
  AO22X1_LVT U2801 ( .A1(n3410), .A2(n3494), .A3(n3409), .A4(\regs[18][22] ), 
        .Y(n1977) );
  AO22X1_LVT U2802 ( .A1(n3410), .A2(wdata[21]), .A3(n3409), .A4(
        \regs[18][21] ), .Y(n1976) );
  AO22X1_LVT U2803 ( .A1(n3412), .A2(n3483), .A3(n3411), .A4(\regs[18][20] ), 
        .Y(n1975) );
  AO22X1_LVT U2804 ( .A1(n3410), .A2(n3496), .A3(n3409), .A4(\regs[18][19] ), 
        .Y(n1974) );
  AO22X1_LVT U2805 ( .A1(n3412), .A2(n3491), .A3(n3411), .A4(\regs[18][18] ), 
        .Y(n1973) );
  AO22X1_LVT U2806 ( .A1(n3410), .A2(wdata[17]), .A3(n3409), .A4(
        \regs[18][17] ), .Y(n1972) );
  AO22X1_LVT U2808 ( .A1(n3410), .A2(wdata[16]), .A3(n3409), .A4(
        \regs[18][16] ), .Y(n1971) );
  AO22X1_LVT U2809 ( .A1(n3410), .A2(n3495), .A3(n3409), .A4(\regs[18][15] ), 
        .Y(n1970) );
  AO22X1_LVT U2810 ( .A1(n3410), .A2(n3498), .A3(n3409), .A4(\regs[18][14] ), 
        .Y(n1969) );
  AO22X1_LVT U2811 ( .A1(n3412), .A2(n3502), .A3(n3411), .A4(\regs[18][13] ), 
        .Y(n1968) );
  AO22X1_LVT U2812 ( .A1(n3412), .A2(wdata[12]), .A3(n3411), .A4(
        \regs[18][12] ), .Y(n1967) );
  AO22X1_LVT U2813 ( .A1(n3410), .A2(wdata[11]), .A3(n3409), .A4(
        \regs[18][11] ), .Y(n1966) );
  AO22X1_LVT U2814 ( .A1(n3412), .A2(n3499), .A3(n3411), .A4(\regs[18][10] ), 
        .Y(n1965) );
  AO22X1_LVT U2815 ( .A1(n3412), .A2(wdata[9]), .A3(n3411), .A4(\regs[18][9] ), 
        .Y(n1964) );
  AO22X1_LVT U2817 ( .A1(n3410), .A2(wdata[8]), .A3(n3409), .A4(\regs[18][8] ), 
        .Y(n1963) );
  AO22X1_LVT U2818 ( .A1(n3410), .A2(wdata[7]), .A3(n3409), .A4(\regs[18][7] ), 
        .Y(n1962) );
  AO22X1_LVT U2819 ( .A1(n3410), .A2(wdata[6]), .A3(n3409), .A4(\regs[18][6] ), 
        .Y(n1961) );
  AO22X1_LVT U2820 ( .A1(n3410), .A2(wdata[5]), .A3(n3409), .A4(\regs[18][5] ), 
        .Y(n1960) );
  AO22X1_LVT U2821 ( .A1(n3410), .A2(wdata[4]), .A3(n3409), .A4(\regs[18][4] ), 
        .Y(n1959) );
  AO22X1_LVT U2822 ( .A1(n3412), .A2(wdata[3]), .A3(n3411), .A4(\regs[18][3] ), 
        .Y(n1958) );
  AO22X1_LVT U2823 ( .A1(n3412), .A2(wdata[2]), .A3(n3411), .A4(\regs[18][2] ), 
        .Y(n1957) );
  AO22X1_LVT U2825 ( .A1(n3412), .A2(wdata[1]), .A3(n3411), .A4(\regs[18][1] ), 
        .Y(n1956) );
  AO22X1_LVT U2826 ( .A1(n3412), .A2(wdata[0]), .A3(n3411), .A4(\regs[18][0] ), 
        .Y(n1955) );
  AO22X1_LVT U2832 ( .A1(n3406), .A2(n3486), .A3(n3405), .A4(\regs[19][31] ), 
        .Y(n1954) );
  AO22X1_LVT U2833 ( .A1(n3404), .A2(wdata[30]), .A3(n3403), .A4(
        \regs[19][30] ), .Y(n1953) );
  AO22X1_LVT U2834 ( .A1(n3404), .A2(n3501), .A3(n3403), .A4(\regs[19][29] ), 
        .Y(n1952) );
  AO22X1_LVT U2835 ( .A1(n3404), .A2(n3500), .A3(n3403), .A4(\regs[19][28] ), 
        .Y(n1951) );
  AO22X1_LVT U2836 ( .A1(n3406), .A2(wdata[27]), .A3(n3405), .A4(
        \regs[19][27] ), .Y(n1950) );
  AO22X1_LVT U2837 ( .A1(n3404), .A2(n3503), .A3(n3403), .A4(\regs[19][26] ), 
        .Y(n1949) );
  AO22X1_LVT U2838 ( .A1(n3406), .A2(wdata[25]), .A3(n3405), .A4(
        \regs[19][25] ), .Y(n1948) );
  AO22X1_LVT U2840 ( .A1(n3408), .A2(n3493), .A3(n3407), .A4(\regs[19][24] ), 
        .Y(n1947) );
  AO22X1_LVT U2841 ( .A1(n3406), .A2(n3497), .A3(n3405), .A4(\regs[19][23] ), 
        .Y(n1946) );
  AO22X1_LVT U2842 ( .A1(n3406), .A2(n3494), .A3(n3405), .A4(\regs[19][22] ), 
        .Y(n1945) );
  AO22X1_LVT U2843 ( .A1(n3408), .A2(wdata[21]), .A3(n3407), .A4(
        \regs[19][21] ), .Y(n1944) );
  AO22X1_LVT U2844 ( .A1(n3406), .A2(n3483), .A3(n3405), .A4(\regs[19][20] ), 
        .Y(n1943) );
  AO22X1_LVT U2845 ( .A1(n3406), .A2(n3496), .A3(n3405), .A4(\regs[19][19] ), 
        .Y(n1942) );
  AO22X1_LVT U2846 ( .A1(n3406), .A2(n3491), .A3(n3405), .A4(\regs[19][18] ), 
        .Y(n1941) );
  AO22X1_LVT U2847 ( .A1(n3408), .A2(wdata[17]), .A3(n3407), .A4(
        \regs[19][17] ), .Y(n1940) );
  AO22X1_LVT U2849 ( .A1(n3404), .A2(wdata[16]), .A3(n3403), .A4(
        \regs[19][16] ), .Y(n1939) );
  AO22X1_LVT U2850 ( .A1(n3404), .A2(n3495), .A3(n3403), .A4(\regs[19][15] ), 
        .Y(n1938) );
  AO22X1_LVT U2851 ( .A1(n3404), .A2(wdata[14]), .A3(n3403), .A4(
        \regs[19][14] ), .Y(n1937) );
  AO22X1_LVT U2852 ( .A1(n3404), .A2(n3502), .A3(n3403), .A4(\regs[19][13] ), 
        .Y(n1936) );
  AO22X1_LVT U2853 ( .A1(n3404), .A2(wdata[12]), .A3(n3403), .A4(
        \regs[19][12] ), .Y(n1935) );
  AO22X1_LVT U2854 ( .A1(n3404), .A2(wdata[11]), .A3(n3403), .A4(
        \regs[19][11] ), .Y(n1934) );
  AO22X1_LVT U2855 ( .A1(n3404), .A2(n3499), .A3(n3403), .A4(\regs[19][10] ), 
        .Y(n1933) );
  AO22X1_LVT U2856 ( .A1(n3404), .A2(wdata[9]), .A3(n3403), .A4(\regs[19][9] ), 
        .Y(n1932) );
  AO22X1_LVT U2858 ( .A1(n3408), .A2(wdata[8]), .A3(n3407), .A4(\regs[19][8] ), 
        .Y(n1931) );
  AO22X1_LVT U2859 ( .A1(n3408), .A2(wdata[7]), .A3(n3407), .A4(\regs[19][7] ), 
        .Y(n1930) );
  AO22X1_LVT U2860 ( .A1(n3408), .A2(wdata[6]), .A3(n3407), .A4(\regs[19][6] ), 
        .Y(n1929) );
  AO22X1_LVT U2861 ( .A1(n3408), .A2(wdata[5]), .A3(n3407), .A4(\regs[19][5] ), 
        .Y(n1928) );
  AO22X1_LVT U2862 ( .A1(n3408), .A2(wdata[4]), .A3(n3407), .A4(\regs[19][4] ), 
        .Y(n1927) );
  AO22X1_LVT U2863 ( .A1(n3408), .A2(wdata[3]), .A3(n3407), .A4(\regs[19][3] ), 
        .Y(n1926) );
  AO22X1_LVT U2864 ( .A1(n3408), .A2(wdata[2]), .A3(n3407), .A4(\regs[19][2] ), 
        .Y(n1925) );
  AO22X1_LVT U2866 ( .A1(n3408), .A2(wdata[1]), .A3(n3407), .A4(\regs[19][1] ), 
        .Y(n1924) );
  AO22X1_LVT U2867 ( .A1(n3408), .A2(wdata[0]), .A3(n3407), .A4(\regs[19][0] ), 
        .Y(n1923) );
  NAND4X0_LVT U2868 ( .A1(n3470), .A2(n3142), .A3(n3192), .A4(n3191), .Y(n3115) );
  AO22X1_LVT U2873 ( .A1(n3308), .A2(n3486), .A3(n3307), .A4(\regs[20][31] ), 
        .Y(n1922) );
  AO22X1_LVT U2874 ( .A1(n3310), .A2(wdata[30]), .A3(n3309), .A4(
        \regs[20][30] ), .Y(n1921) );
  AO22X1_LVT U2875 ( .A1(n3310), .A2(n3501), .A3(n3309), .A4(\regs[20][29] ), 
        .Y(n1920) );
  AO22X1_LVT U2876 ( .A1(n3308), .A2(n3500), .A3(n3307), .A4(\regs[20][28] ), 
        .Y(n1919) );
  AO22X1_LVT U2877 ( .A1(n3308), .A2(wdata[27]), .A3(n3307), .A4(
        \regs[20][27] ), .Y(n1918) );
  AO22X1_LVT U2878 ( .A1(n3310), .A2(n3503), .A3(n3309), .A4(\regs[20][26] ), 
        .Y(n1917) );
  AO22X1_LVT U2879 ( .A1(n3308), .A2(wdata[25]), .A3(n3307), .A4(
        \regs[20][25] ), .Y(n1916) );
  AO22X1_LVT U2881 ( .A1(n3310), .A2(n3493), .A3(n3309), .A4(\regs[20][24] ), 
        .Y(n1915) );
  AO22X1_LVT U2882 ( .A1(n3308), .A2(n3497), .A3(n3307), .A4(\regs[20][23] ), 
        .Y(n1914) );
  AO22X1_LVT U2883 ( .A1(n3308), .A2(n3494), .A3(n3307), .A4(\regs[20][22] ), 
        .Y(n1913) );
  AO22X1_LVT U2884 ( .A1(n3308), .A2(wdata[21]), .A3(n3307), .A4(
        \regs[20][21] ), .Y(n1912) );
  AO22X1_LVT U2885 ( .A1(n3308), .A2(n3483), .A3(n3307), .A4(\regs[20][20] ), 
        .Y(n1911) );
  AO22X1_LVT U2886 ( .A1(n3310), .A2(n3496), .A3(n3309), .A4(\regs[20][19] ), 
        .Y(n1910) );
  AO22X1_LVT U2887 ( .A1(n3310), .A2(n3491), .A3(n3309), .A4(\regs[20][18] ), 
        .Y(n1909) );
  AO22X1_LVT U2888 ( .A1(n3310), .A2(wdata[17]), .A3(n3309), .A4(
        \regs[20][17] ), .Y(n1908) );
  AO22X1_LVT U2890 ( .A1(n3308), .A2(wdata[16]), .A3(n3307), .A4(
        \regs[20][16] ), .Y(n1907) );
  AO22X1_LVT U2891 ( .A1(n3310), .A2(n3495), .A3(n3309), .A4(\regs[20][15] ), 
        .Y(n1906) );
  AO22X1_LVT U2892 ( .A1(n3308), .A2(n3498), .A3(n3307), .A4(\regs[20][14] ), 
        .Y(n1905) );
  AO22X1_LVT U2893 ( .A1(n3308), .A2(n3502), .A3(n3307), .A4(\regs[20][13] ), 
        .Y(n1904) );
  AO22X1_LVT U2894 ( .A1(n3310), .A2(wdata[12]), .A3(n3309), .A4(
        \regs[20][12] ), .Y(n1903) );
  AO22X1_LVT U2895 ( .A1(n3308), .A2(wdata[11]), .A3(n3307), .A4(
        \regs[20][11] ), .Y(n1902) );
  AO22X1_LVT U2896 ( .A1(n3308), .A2(n3499), .A3(n3307), .A4(\regs[20][10] ), 
        .Y(n1901) );
  AO22X1_LVT U2897 ( .A1(n3310), .A2(wdata[9]), .A3(n3309), .A4(\regs[20][9] ), 
        .Y(n1900) );
  AO22X1_LVT U2899 ( .A1(n3310), .A2(wdata[8]), .A3(n3309), .A4(\regs[20][8] ), 
        .Y(n1899) );
  AO22X1_LVT U2900 ( .A1(n3310), .A2(wdata[7]), .A3(n3309), .A4(\regs[20][7] ), 
        .Y(n1898) );
  AO22X1_LVT U2901 ( .A1(n3310), .A2(wdata[6]), .A3(n3309), .A4(\regs[20][6] ), 
        .Y(n1897) );
  AO22X1_LVT U2902 ( .A1(n3310), .A2(wdata[5]), .A3(n3309), .A4(\regs[20][5] ), 
        .Y(n1896) );
  AO22X1_LVT U2903 ( .A1(n3310), .A2(wdata[4]), .A3(n3309), .A4(\regs[20][4] ), 
        .Y(n1895) );
  AO22X1_LVT U2904 ( .A1(n3310), .A2(wdata[3]), .A3(n3309), .A4(\regs[20][3] ), 
        .Y(n1894) );
  AO22X1_LVT U2905 ( .A1(n3310), .A2(wdata[2]), .A3(n3309), .A4(\regs[20][2] ), 
        .Y(n1893) );
  AO22X1_LVT U2907 ( .A1(n3310), .A2(wdata[1]), .A3(n3309), .A4(\regs[20][1] ), 
        .Y(n1892) );
  AO22X1_LVT U2908 ( .A1(n3310), .A2(wdata[0]), .A3(n3309), .A4(\regs[20][0] ), 
        .Y(n1891) );
  AO22X1_LVT U2914 ( .A1(n3344), .A2(wdata[31]), .A3(n3343), .A4(
        \regs[21][31] ), .Y(n1890) );
  AO22X1_LVT U2915 ( .A1(n3344), .A2(wdata[30]), .A3(n3343), .A4(
        \regs[21][30] ), .Y(n1889) );
  AO22X1_LVT U2916 ( .A1(n3344), .A2(n3501), .A3(n3343), .A4(\regs[21][29] ), 
        .Y(n1888) );
  AO22X1_LVT U2917 ( .A1(n3344), .A2(n3500), .A3(n3343), .A4(\regs[21][28] ), 
        .Y(n1887) );
  AO22X1_LVT U2918 ( .A1(n3344), .A2(wdata[27]), .A3(n3343), .A4(
        \regs[21][27] ), .Y(n1886) );
  AO22X1_LVT U2919 ( .A1(n3344), .A2(n3503), .A3(n3343), .A4(\regs[21][26] ), 
        .Y(n1885) );
  AO22X1_LVT U2920 ( .A1(n3344), .A2(wdata[25]), .A3(n3343), .A4(
        \regs[21][25] ), .Y(n1884) );
  AO22X1_LVT U2922 ( .A1(n3346), .A2(n3493), .A3(n3345), .A4(\regs[21][24] ), 
        .Y(n1883) );
  AO22X1_LVT U2923 ( .A1(n3344), .A2(n3497), .A3(n3343), .A4(\regs[21][23] ), 
        .Y(n1882) );
  AO22X1_LVT U2924 ( .A1(n3346), .A2(n3494), .A3(n3345), .A4(\regs[21][22] ), 
        .Y(n1881) );
  AO22X1_LVT U2925 ( .A1(n3346), .A2(wdata[21]), .A3(n3345), .A4(
        \regs[21][21] ), .Y(n1880) );
  AO22X1_LVT U2926 ( .A1(n3344), .A2(n3492), .A3(n3343), .A4(\regs[21][20] ), 
        .Y(n1879) );
  AO22X1_LVT U2927 ( .A1(n3344), .A2(n3496), .A3(n3343), .A4(\regs[21][19] ), 
        .Y(n1878) );
  AO22X1_LVT U2928 ( .A1(n3346), .A2(n3491), .A3(n3345), .A4(\regs[21][18] ), 
        .Y(n1877) );
  AO22X1_LVT U2929 ( .A1(n3346), .A2(wdata[17]), .A3(n3345), .A4(
        \regs[21][17] ), .Y(n1876) );
  AO22X1_LVT U2931 ( .A1(n3344), .A2(wdata[16]), .A3(n3343), .A4(
        \regs[21][16] ), .Y(n1875) );
  AO22X1_LVT U2932 ( .A1(n3344), .A2(n3495), .A3(n3343), .A4(\regs[21][15] ), 
        .Y(n1874) );
  AO22X1_LVT U2933 ( .A1(n3344), .A2(n3498), .A3(n3343), .A4(\regs[21][14] ), 
        .Y(n1873) );
  AO22X1_LVT U2934 ( .A1(n3344), .A2(n3502), .A3(n3343), .A4(\regs[21][13] ), 
        .Y(n1872) );
  AO22X1_LVT U2935 ( .A1(n3344), .A2(wdata[12]), .A3(n3343), .A4(
        \regs[21][12] ), .Y(n1871) );
  AO22X1_LVT U2936 ( .A1(n3344), .A2(wdata[11]), .A3(n3343), .A4(
        \regs[21][11] ), .Y(n1870) );
  AO22X1_LVT U2937 ( .A1(n3344), .A2(n3499), .A3(n3343), .A4(\regs[21][10] ), 
        .Y(n1869) );
  AO22X1_LVT U2938 ( .A1(n3344), .A2(wdata[9]), .A3(n3343), .A4(\regs[21][9] ), 
        .Y(n1868) );
  AO22X1_LVT U2940 ( .A1(n3346), .A2(wdata[8]), .A3(n3345), .A4(\regs[21][8] ), 
        .Y(n1867) );
  AO22X1_LVT U2941 ( .A1(n3346), .A2(wdata[7]), .A3(n3345), .A4(\regs[21][7] ), 
        .Y(n1866) );
  AO22X1_LVT U2942 ( .A1(n3346), .A2(wdata[6]), .A3(n3345), .A4(\regs[21][6] ), 
        .Y(n1865) );
  AO22X1_LVT U2943 ( .A1(n3346), .A2(wdata[5]), .A3(n3345), .A4(\regs[21][5] ), 
        .Y(n1864) );
  AO22X1_LVT U2944 ( .A1(n3346), .A2(wdata[4]), .A3(n3345), .A4(\regs[21][4] ), 
        .Y(n1863) );
  AO22X1_LVT U2945 ( .A1(n3346), .A2(wdata[3]), .A3(n3345), .A4(\regs[21][3] ), 
        .Y(n1862) );
  AO22X1_LVT U2946 ( .A1(n3346), .A2(wdata[2]), .A3(n3345), .A4(\regs[21][2] ), 
        .Y(n1861) );
  AO22X1_LVT U2948 ( .A1(n3346), .A2(wdata[1]), .A3(n3345), .A4(\regs[21][1] ), 
        .Y(n1860) );
  AO22X1_LVT U2949 ( .A1(n3346), .A2(wdata[0]), .A3(n3345), .A4(\regs[21][0] ), 
        .Y(n1859) );
  NAND3X0_LVT U2950 ( .A1(n3470), .A2(n3212), .A3(n3142), .Y(n3133) );
  AO22X1_LVT U2955 ( .A1(n3340), .A2(n3486), .A3(n3339), .A4(\regs[22][31] ), 
        .Y(n1858) );
  AO22X1_LVT U2956 ( .A1(n3342), .A2(wdata[30]), .A3(n3341), .A4(
        \regs[22][30] ), .Y(n1857) );
  AO22X1_LVT U2957 ( .A1(n3342), .A2(n3501), .A3(n3341), .A4(\regs[22][29] ), 
        .Y(n1856) );
  AO22X1_LVT U2958 ( .A1(n3342), .A2(n3500), .A3(n3341), .A4(\regs[22][28] ), 
        .Y(n1855) );
  AO22X1_LVT U2959 ( .A1(n3342), .A2(wdata[27]), .A3(n3341), .A4(
        \regs[22][27] ), .Y(n1854) );
  AO22X1_LVT U2960 ( .A1(n3342), .A2(n3503), .A3(n3341), .A4(\regs[22][26] ), 
        .Y(n1853) );
  AO22X1_LVT U2961 ( .A1(n3342), .A2(wdata[25]), .A3(n3341), .A4(
        \regs[22][25] ), .Y(n1852) );
  AO22X1_LVT U2963 ( .A1(n3340), .A2(n3493), .A3(n3339), .A4(\regs[22][24] ), 
        .Y(n1851) );
  AO22X1_LVT U2964 ( .A1(n3340), .A2(n3497), .A3(n3339), .A4(\regs[22][23] ), 
        .Y(n1850) );
  AO22X1_LVT U2965 ( .A1(n3340), .A2(n3494), .A3(n3339), .A4(\regs[22][22] ), 
        .Y(n1849) );
  AO22X1_LVT U2966 ( .A1(n3340), .A2(wdata[21]), .A3(n3339), .A4(
        \regs[22][21] ), .Y(n1848) );
  AO22X1_LVT U2967 ( .A1(n3340), .A2(n3483), .A3(n3339), .A4(\regs[22][20] ), 
        .Y(n1847) );
  AO22X1_LVT U2968 ( .A1(n3340), .A2(n3496), .A3(n3339), .A4(\regs[22][19] ), 
        .Y(n1846) );
  AO22X1_LVT U2969 ( .A1(n3340), .A2(n3491), .A3(n3339), .A4(\regs[22][18] ), 
        .Y(n1845) );
  AO22X1_LVT U2970 ( .A1(n3340), .A2(wdata[17]), .A3(n3339), .A4(
        \regs[22][17] ), .Y(n1844) );
  AO22X1_LVT U2972 ( .A1(n3342), .A2(wdata[16]), .A3(n3341), .A4(
        \regs[22][16] ), .Y(n1843) );
  AO22X1_LVT U2973 ( .A1(n3340), .A2(n3495), .A3(n3339), .A4(\regs[22][15] ), 
        .Y(n1842) );
  AO22X1_LVT U2974 ( .A1(n3340), .A2(n3498), .A3(n3339), .A4(\regs[22][14] ), 
        .Y(n1841) );
  AO22X1_LVT U2975 ( .A1(n3342), .A2(n3502), .A3(n3341), .A4(\regs[22][13] ), 
        .Y(n1840) );
  AO22X1_LVT U2976 ( .A1(n3342), .A2(wdata[12]), .A3(n3341), .A4(
        \regs[22][12] ), .Y(n1839) );
  AO22X1_LVT U2977 ( .A1(n3340), .A2(wdata[11]), .A3(n3339), .A4(
        \regs[22][11] ), .Y(n1838) );
  AO22X1_LVT U2978 ( .A1(n3342), .A2(n3499), .A3(n3341), .A4(\regs[22][10] ), 
        .Y(n1837) );
  AO22X1_LVT U2979 ( .A1(n3340), .A2(wdata[9]), .A3(n3339), .A4(\regs[22][9] ), 
        .Y(n1836) );
  AO22X1_LVT U2981 ( .A1(n3342), .A2(wdata[8]), .A3(n3341), .A4(\regs[22][8] ), 
        .Y(n1835) );
  AO22X1_LVT U2982 ( .A1(n3340), .A2(wdata[7]), .A3(n3339), .A4(\regs[22][7] ), 
        .Y(n1834) );
  AO22X1_LVT U2983 ( .A1(n3340), .A2(wdata[6]), .A3(n3339), .A4(\regs[22][6] ), 
        .Y(n1833) );
  AO22X1_LVT U2984 ( .A1(n3340), .A2(wdata[5]), .A3(n3339), .A4(\regs[22][5] ), 
        .Y(n1832) );
  AO22X1_LVT U2985 ( .A1(n3340), .A2(wdata[4]), .A3(n3339), .A4(\regs[22][4] ), 
        .Y(n1831) );
  AO22X1_LVT U2986 ( .A1(n3342), .A2(wdata[3]), .A3(n3341), .A4(\regs[22][3] ), 
        .Y(n1830) );
  AO22X1_LVT U2987 ( .A1(n3340), .A2(wdata[2]), .A3(n3339), .A4(\regs[22][2] ), 
        .Y(n1829) );
  AO22X1_LVT U2989 ( .A1(n3340), .A2(wdata[1]), .A3(n3339), .A4(\regs[22][1] ), 
        .Y(n1828) );
  AO22X1_LVT U2990 ( .A1(n3340), .A2(wdata[0]), .A3(n3339), .A4(\regs[22][0] ), 
        .Y(n1827) );
  AO22X1_LVT U2996 ( .A1(n3334), .A2(n3486), .A3(n3333), .A4(\regs[23][31] ), 
        .Y(n1826) );
  AO22X1_LVT U2997 ( .A1(n3334), .A2(wdata[30]), .A3(n3333), .A4(
        \regs[23][30] ), .Y(n1825) );
  AO22X1_LVT U2998 ( .A1(n3334), .A2(n3501), .A3(n3333), .A4(\regs[23][29] ), 
        .Y(n1824) );
  AO22X1_LVT U2999 ( .A1(n3334), .A2(n3500), .A3(n3333), .A4(\regs[23][28] ), 
        .Y(n1823) );
  AO22X1_LVT U3000 ( .A1(n3334), .A2(wdata[27]), .A3(n3333), .A4(
        \regs[23][27] ), .Y(n1822) );
  AO22X1_LVT U3001 ( .A1(n3334), .A2(n3503), .A3(n3333), .A4(\regs[23][26] ), 
        .Y(n1821) );
  AO22X1_LVT U3002 ( .A1(n3334), .A2(wdata[25]), .A3(n3333), .A4(
        \regs[23][25] ), .Y(n1820) );
  AO22X1_LVT U3004 ( .A1(n3336), .A2(n3493), .A3(n3335), .A4(\regs[23][24] ), 
        .Y(n1819) );
  AO22X1_LVT U3005 ( .A1(n3336), .A2(n3497), .A3(n3335), .A4(\regs[23][23] ), 
        .Y(n1818) );
  AO22X1_LVT U3006 ( .A1(n3336), .A2(n3494), .A3(n3335), .A4(\regs[23][22] ), 
        .Y(n1817) );
  AO22X1_LVT U3007 ( .A1(n3336), .A2(wdata[21]), .A3(n3335), .A4(
        \regs[23][21] ), .Y(n1816) );
  AO22X1_LVT U3008 ( .A1(n3336), .A2(n3483), .A3(n3335), .A4(\regs[23][20] ), 
        .Y(n1815) );
  AO22X1_LVT U3009 ( .A1(n3336), .A2(n3496), .A3(n3335), .A4(\regs[23][19] ), 
        .Y(n1814) );
  AO22X1_LVT U3010 ( .A1(n3336), .A2(n3491), .A3(n3335), .A4(\regs[23][18] ), 
        .Y(n1813) );
  AO22X1_LVT U3011 ( .A1(n3336), .A2(wdata[17]), .A3(n3335), .A4(
        \regs[23][17] ), .Y(n1812) );
  AO22X1_LVT U3013 ( .A1(n3334), .A2(wdata[16]), .A3(n3333), .A4(
        \regs[23][16] ), .Y(n1811) );
  AO22X1_LVT U3014 ( .A1(n3334), .A2(n3495), .A3(n3333), .A4(\regs[23][15] ), 
        .Y(n1810) );
  AO22X1_LVT U3015 ( .A1(n3334), .A2(n3498), .A3(n3333), .A4(\regs[23][14] ), 
        .Y(n1809) );
  AO22X1_LVT U3016 ( .A1(n3334), .A2(n3502), .A3(n3333), .A4(\regs[23][13] ), 
        .Y(n1808) );
  AO22X1_LVT U3017 ( .A1(n3334), .A2(wdata[12]), .A3(n3333), .A4(
        \regs[23][12] ), .Y(n1807) );
  AO22X1_LVT U3018 ( .A1(n3334), .A2(wdata[11]), .A3(n3333), .A4(
        \regs[23][11] ), .Y(n1806) );
  AO22X1_LVT U3019 ( .A1(n3334), .A2(n3499), .A3(n3333), .A4(\regs[23][10] ), 
        .Y(n1805) );
  AO22X1_LVT U3020 ( .A1(n3334), .A2(wdata[9]), .A3(n3333), .A4(\regs[23][9] ), 
        .Y(n1804) );
  AO22X1_LVT U3022 ( .A1(n3338), .A2(wdata[8]), .A3(n3337), .A4(\regs[23][8] ), 
        .Y(n1803) );
  AO22X1_LVT U3023 ( .A1(n3338), .A2(wdata[7]), .A3(n3337), .A4(\regs[23][7] ), 
        .Y(n1802) );
  AO22X1_LVT U3024 ( .A1(n3338), .A2(wdata[6]), .A3(n3337), .A4(\regs[23][6] ), 
        .Y(n1801) );
  AO22X1_LVT U3025 ( .A1(n3338), .A2(wdata[5]), .A3(n3337), .A4(\regs[23][5] ), 
        .Y(n1800) );
  AO22X1_LVT U3026 ( .A1(n3338), .A2(wdata[4]), .A3(n3337), .A4(\regs[23][4] ), 
        .Y(n1799) );
  AO22X1_LVT U3027 ( .A1(n3338), .A2(wdata[3]), .A3(n3337), .A4(\regs[23][3] ), 
        .Y(n1798) );
  AO22X1_LVT U3028 ( .A1(n3338), .A2(wdata[2]), .A3(n3337), .A4(\regs[23][2] ), 
        .Y(n1797) );
  AO22X1_LVT U3030 ( .A1(n3336), .A2(wdata[1]), .A3(n3335), .A4(\regs[23][1] ), 
        .Y(n1796) );
  AO22X1_LVT U3031 ( .A1(n3336), .A2(wdata[0]), .A3(n3335), .A4(\regs[23][0] ), 
        .Y(n1795) );
  AND4X1_LVT U3032 ( .A1(waddr[4]), .A2(waddr[3]), .A3(we), .A4(n3297), .Y(
        n3254) );
  AND2X1_LVT U3033 ( .A1(n3254), .A2(n3298), .Y(n3181) );
  AO22X1_LVT U3039 ( .A1(n3330), .A2(wdata[31]), .A3(n3329), .A4(
        \regs[24][31] ), .Y(n1794) );
  AO22X1_LVT U3040 ( .A1(n3330), .A2(wdata[30]), .A3(n3329), .A4(
        \regs[24][30] ), .Y(n1793) );
  AO22X1_LVT U3041 ( .A1(n3330), .A2(n3501), .A3(n3329), .A4(\regs[24][29] ), 
        .Y(n1792) );
  AO22X1_LVT U3042 ( .A1(n3330), .A2(n3500), .A3(n3329), .A4(\regs[24][28] ), 
        .Y(n1791) );
  AO22X1_LVT U3043 ( .A1(n3330), .A2(wdata[27]), .A3(n3329), .A4(
        \regs[24][27] ), .Y(n1790) );
  AO22X1_LVT U3044 ( .A1(n3330), .A2(n3503), .A3(n3329), .A4(\regs[24][26] ), 
        .Y(n1789) );
  AO22X1_LVT U3045 ( .A1(n3330), .A2(wdata[25]), .A3(n3329), .A4(
        \regs[24][25] ), .Y(n1788) );
  AO22X1_LVT U3047 ( .A1(n3332), .A2(n3493), .A3(n3331), .A4(\regs[24][24] ), 
        .Y(n1787) );
  AO22X1_LVT U3048 ( .A1(n3332), .A2(n3497), .A3(n3331), .A4(\regs[24][23] ), 
        .Y(n1786) );
  AO22X1_LVT U3049 ( .A1(n3332), .A2(n3494), .A3(n3331), .A4(\regs[24][22] ), 
        .Y(n1785) );
  AO22X1_LVT U3050 ( .A1(n3332), .A2(wdata[21]), .A3(n3331), .A4(
        \regs[24][21] ), .Y(n1784) );
  AO22X1_LVT U3051 ( .A1(n3332), .A2(n3483), .A3(n3331), .A4(\regs[24][20] ), 
        .Y(n1783) );
  AO22X1_LVT U3052 ( .A1(n3332), .A2(n3496), .A3(n3331), .A4(\regs[24][19] ), 
        .Y(n1782) );
  AO22X1_LVT U3053 ( .A1(n3332), .A2(n3491), .A3(n3331), .A4(\regs[24][18] ), 
        .Y(n1781) );
  AO22X1_LVT U3054 ( .A1(n3332), .A2(wdata[17]), .A3(n3331), .A4(
        \regs[24][17] ), .Y(n1780) );
  AO22X1_LVT U3056 ( .A1(n3330), .A2(wdata[16]), .A3(n3329), .A4(
        \regs[24][16] ), .Y(n1779) );
  AO22X1_LVT U3057 ( .A1(n3330), .A2(n3495), .A3(n3329), .A4(\regs[24][15] ), 
        .Y(n1778) );
  AO22X1_LVT U3058 ( .A1(n3330), .A2(n3498), .A3(n3329), .A4(\regs[24][14] ), 
        .Y(n1777) );
  AO22X1_LVT U3059 ( .A1(n3330), .A2(n3502), .A3(n3329), .A4(\regs[24][13] ), 
        .Y(n1776) );
  AO22X1_LVT U3060 ( .A1(n3330), .A2(wdata[12]), .A3(n3329), .A4(
        \regs[24][12] ), .Y(n1775) );
  AO22X1_LVT U3061 ( .A1(n3330), .A2(wdata[11]), .A3(n3329), .A4(
        \regs[24][11] ), .Y(n1774) );
  AO22X1_LVT U3062 ( .A1(n3330), .A2(n3499), .A3(n3329), .A4(\regs[24][10] ), 
        .Y(n1773) );
  AO22X1_LVT U3063 ( .A1(n3330), .A2(wdata[9]), .A3(n3329), .A4(\regs[24][9] ), 
        .Y(n1772) );
  AO22X1_LVT U3065 ( .A1(n3332), .A2(wdata[8]), .A3(n3331), .A4(\regs[24][8] ), 
        .Y(n1771) );
  AO22X1_LVT U3066 ( .A1(n3332), .A2(wdata[7]), .A3(n3331), .A4(\regs[24][7] ), 
        .Y(n1770) );
  AO22X1_LVT U3067 ( .A1(n3332), .A2(wdata[6]), .A3(n3331), .A4(\regs[24][6] ), 
        .Y(n1769) );
  AO22X1_LVT U3068 ( .A1(n3332), .A2(wdata[5]), .A3(n3331), .A4(\regs[24][5] ), 
        .Y(n1768) );
  AO22X1_LVT U3069 ( .A1(n3332), .A2(wdata[4]), .A3(n3331), .A4(\regs[24][4] ), 
        .Y(n1767) );
  AO22X1_LVT U3070 ( .A1(n3332), .A2(wdata[3]), .A3(n3331), .A4(\regs[24][3] ), 
        .Y(n1766) );
  AO22X1_LVT U3071 ( .A1(n3332), .A2(wdata[2]), .A3(n3331), .A4(\regs[24][2] ), 
        .Y(n1765) );
  AO22X1_LVT U3073 ( .A1(n3332), .A2(wdata[1]), .A3(n3331), .A4(\regs[24][1] ), 
        .Y(n1764) );
  AO22X1_LVT U3074 ( .A1(n3332), .A2(wdata[0]), .A3(n3331), .A4(\regs[24][0] ), 
        .Y(n1763) );
  NAND2X0_LVT U3075 ( .A1(n3202), .A2(n3181), .Y(n3163) );
  AO22X1_LVT U3080 ( .A1(n3390), .A2(n3486), .A3(n3389), .A4(\regs[25][31] ), 
        .Y(n1762) );
  AO22X1_LVT U3081 ( .A1(n3392), .A2(wdata[30]), .A3(n3391), .A4(
        \regs[25][30] ), .Y(n1761) );
  AO22X1_LVT U3082 ( .A1(n3390), .A2(n3501), .A3(n3389), .A4(\regs[25][29] ), 
        .Y(n1760) );
  AO22X1_LVT U3083 ( .A1(n3392), .A2(n3500), .A3(n3391), .A4(\regs[25][28] ), 
        .Y(n1759) );
  AO22X1_LVT U3084 ( .A1(n3392), .A2(wdata[27]), .A3(n3391), .A4(
        \regs[25][27] ), .Y(n1758) );
  AO22X1_LVT U3085 ( .A1(n3392), .A2(n3503), .A3(n3391), .A4(\regs[25][26] ), 
        .Y(n1757) );
  AO22X1_LVT U3086 ( .A1(n3390), .A2(wdata[25]), .A3(n3389), .A4(
        \regs[25][25] ), .Y(n1756) );
  AO22X1_LVT U3088 ( .A1(n3390), .A2(n3493), .A3(n3389), .A4(\regs[25][24] ), 
        .Y(n1755) );
  AO22X1_LVT U3089 ( .A1(n3390), .A2(n3497), .A3(n3389), .A4(\regs[25][23] ), 
        .Y(n1754) );
  AO22X1_LVT U3090 ( .A1(n3390), .A2(n3494), .A3(n3389), .A4(\regs[25][22] ), 
        .Y(n1753) );
  AO22X1_LVT U3091 ( .A1(n3392), .A2(wdata[21]), .A3(n3391), .A4(
        \regs[25][21] ), .Y(n1752) );
  AO22X1_LVT U3092 ( .A1(n3392), .A2(n3483), .A3(n3391), .A4(\regs[25][20] ), 
        .Y(n1751) );
  AO22X1_LVT U3093 ( .A1(n3392), .A2(n3496), .A3(n3391), .A4(\regs[25][19] ), 
        .Y(n1750) );
  AO22X1_LVT U3094 ( .A1(n3390), .A2(n3491), .A3(n3389), .A4(\regs[25][18] ), 
        .Y(n1749) );
  AO22X1_LVT U3095 ( .A1(n3390), .A2(wdata[17]), .A3(n3389), .A4(
        \regs[25][17] ), .Y(n1748) );
  AO22X1_LVT U3097 ( .A1(n3390), .A2(wdata[16]), .A3(n3389), .A4(
        \regs[25][16] ), .Y(n1747) );
  AO22X1_LVT U3098 ( .A1(n3390), .A2(n3495), .A3(n3389), .A4(\regs[25][15] ), 
        .Y(n1746) );
  AO22X1_LVT U3099 ( .A1(n3390), .A2(n3498), .A3(n3389), .A4(\regs[25][14] ), 
        .Y(n1745) );
  AO22X1_LVT U3100 ( .A1(n3390), .A2(n3502), .A3(n3389), .A4(\regs[25][13] ), 
        .Y(n1744) );
  AO22X1_LVT U3101 ( .A1(n3390), .A2(wdata[12]), .A3(n3389), .A4(
        \regs[25][12] ), .Y(n1743) );
  AO22X1_LVT U3102 ( .A1(n3390), .A2(wdata[11]), .A3(n3389), .A4(
        \regs[25][11] ), .Y(n1742) );
  AO22X1_LVT U3103 ( .A1(n3392), .A2(n3499), .A3(n3391), .A4(\regs[25][10] ), 
        .Y(n1741) );
  AO22X1_LVT U3104 ( .A1(n3390), .A2(wdata[9]), .A3(n3389), .A4(\regs[25][9] ), 
        .Y(n1740) );
  AO22X1_LVT U3106 ( .A1(n3392), .A2(wdata[8]), .A3(n3391), .A4(\regs[25][8] ), 
        .Y(n1739) );
  AO22X1_LVT U3107 ( .A1(n3392), .A2(wdata[7]), .A3(n3391), .A4(\regs[25][7] ), 
        .Y(n1738) );
  AO22X1_LVT U3108 ( .A1(n3392), .A2(wdata[6]), .A3(n3391), .A4(\regs[25][6] ), 
        .Y(n1737) );
  AO22X1_LVT U3109 ( .A1(n3392), .A2(wdata[5]), .A3(n3391), .A4(\regs[25][5] ), 
        .Y(n1736) );
  AO22X1_LVT U3110 ( .A1(n3392), .A2(wdata[4]), .A3(n3391), .A4(\regs[25][4] ), 
        .Y(n1735) );
  AO22X1_LVT U3111 ( .A1(n3392), .A2(wdata[3]), .A3(n3391), .A4(\regs[25][3] ), 
        .Y(n1734) );
  AO22X1_LVT U3112 ( .A1(n3392), .A2(wdata[2]), .A3(n3391), .A4(\regs[25][2] ), 
        .Y(n1733) );
  AO22X1_LVT U3114 ( .A1(n3392), .A2(wdata[1]), .A3(n3391), .A4(\regs[25][1] ), 
        .Y(n1732) );
  AO22X1_LVT U3115 ( .A1(n3392), .A2(wdata[0]), .A3(n3391), .A4(\regs[25][0] ), 
        .Y(n1731) );
  NAND2X0_LVT U3116 ( .A1(n3212), .A2(n3181), .Y(n3172) );
  AO22X1_LVT U3121 ( .A1(n3386), .A2(wdata[31]), .A3(n3385), .A4(
        \regs[26][31] ), .Y(n1730) );
  AO22X1_LVT U3122 ( .A1(n3386), .A2(wdata[30]), .A3(n3385), .A4(
        \regs[26][30] ), .Y(n1729) );
  AO22X1_LVT U3123 ( .A1(n3386), .A2(n3501), .A3(n3385), .A4(\regs[26][29] ), 
        .Y(n1728) );
  AO22X1_LVT U3124 ( .A1(n3386), .A2(n3500), .A3(n3385), .A4(\regs[26][28] ), 
        .Y(n1727) );
  AO22X1_LVT U3125 ( .A1(n3386), .A2(wdata[27]), .A3(n3385), .A4(
        \regs[26][27] ), .Y(n1726) );
  AO22X1_LVT U3126 ( .A1(n3386), .A2(n3503), .A3(n3385), .A4(\regs[26][26] ), 
        .Y(n1725) );
  AO22X1_LVT U3127 ( .A1(n3386), .A2(wdata[25]), .A3(n3385), .A4(
        \regs[26][25] ), .Y(n1724) );
  AO22X1_LVT U3129 ( .A1(n3388), .A2(n3493), .A3(n3387), .A4(\regs[26][24] ), 
        .Y(n1723) );
  AO22X1_LVT U3130 ( .A1(n3386), .A2(n3497), .A3(n3385), .A4(\regs[26][23] ), 
        .Y(n1722) );
  AO22X1_LVT U3131 ( .A1(n3386), .A2(n3494), .A3(n3385), .A4(\regs[26][22] ), 
        .Y(n1721) );
  AO22X1_LVT U3132 ( .A1(n3388), .A2(wdata[21]), .A3(n3387), .A4(
        \regs[26][21] ), .Y(n1720) );
  AO22X1_LVT U3133 ( .A1(n3388), .A2(n3492), .A3(n3387), .A4(\regs[26][20] ), 
        .Y(n1719) );
  AO22X1_LVT U3134 ( .A1(n3386), .A2(n3496), .A3(n3385), .A4(\regs[26][19] ), 
        .Y(n1718) );
  AO22X1_LVT U3135 ( .A1(n3386), .A2(n3491), .A3(n3385), .A4(\regs[26][18] ), 
        .Y(n1717) );
  AO22X1_LVT U3136 ( .A1(n3388), .A2(wdata[17]), .A3(n3387), .A4(
        \regs[26][17] ), .Y(n1716) );
  AO22X1_LVT U3138 ( .A1(n3386), .A2(wdata[16]), .A3(n3385), .A4(
        \regs[26][16] ), .Y(n1715) );
  AO22X1_LVT U3139 ( .A1(n3386), .A2(n3495), .A3(n3385), .A4(\regs[26][15] ), 
        .Y(n1714) );
  AO22X1_LVT U3140 ( .A1(n3386), .A2(n3498), .A3(n3385), .A4(\regs[26][14] ), 
        .Y(n1713) );
  AO22X1_LVT U3141 ( .A1(n3386), .A2(n3502), .A3(n3385), .A4(\regs[26][13] ), 
        .Y(n1712) );
  AO22X1_LVT U3142 ( .A1(n3386), .A2(wdata[12]), .A3(n3385), .A4(
        \regs[26][12] ), .Y(n1711) );
  AO22X1_LVT U3143 ( .A1(n3386), .A2(wdata[11]), .A3(n3385), .A4(
        \regs[26][11] ), .Y(n1710) );
  AO22X1_LVT U3144 ( .A1(n3386), .A2(n3499), .A3(n3385), .A4(\regs[26][10] ), 
        .Y(n1709) );
  AO22X1_LVT U3145 ( .A1(n3386), .A2(wdata[9]), .A3(n3385), .A4(\regs[26][9] ), 
        .Y(n1708) );
  AO22X1_LVT U3147 ( .A1(n3388), .A2(wdata[8]), .A3(n3387), .A4(\regs[26][8] ), 
        .Y(n1707) );
  AO22X1_LVT U3148 ( .A1(n3388), .A2(wdata[7]), .A3(n3387), .A4(\regs[26][7] ), 
        .Y(n1706) );
  AO22X1_LVT U3149 ( .A1(n3388), .A2(wdata[6]), .A3(n3387), .A4(\regs[26][6] ), 
        .Y(n1705) );
  AO22X1_LVT U3150 ( .A1(n3388), .A2(wdata[5]), .A3(n3387), .A4(\regs[26][5] ), 
        .Y(n1704) );
  AO22X1_LVT U3151 ( .A1(n3388), .A2(wdata[4]), .A3(n3387), .A4(\regs[26][4] ), 
        .Y(n1703) );
  AO22X1_LVT U3152 ( .A1(n3388), .A2(wdata[3]), .A3(n3387), .A4(\regs[26][3] ), 
        .Y(n1702) );
  AO22X1_LVT U3153 ( .A1(n3388), .A2(wdata[2]), .A3(n3387), .A4(\regs[26][2] ), 
        .Y(n1701) );
  AO22X1_LVT U3155 ( .A1(n3388), .A2(wdata[1]), .A3(n3387), .A4(\regs[26][1] ), 
        .Y(n1700) );
  AO22X1_LVT U3156 ( .A1(n3388), .A2(wdata[0]), .A3(n3387), .A4(\regs[26][0] ), 
        .Y(n1699) );
  AO22X1_LVT U3162 ( .A1(n3384), .A2(n3486), .A3(n3383), .A4(\regs[27][31] ), 
        .Y(n1698) );
  AO22X1_LVT U3163 ( .A1(n3380), .A2(wdata[30]), .A3(n3379), .A4(
        \regs[27][30] ), .Y(n1697) );
  AO22X1_LVT U3164 ( .A1(n3380), .A2(n3501), .A3(n3379), .A4(\regs[27][29] ), 
        .Y(n1696) );
  AO22X1_LVT U3165 ( .A1(n3380), .A2(n3500), .A3(n3379), .A4(\regs[27][28] ), 
        .Y(n1695) );
  AO22X1_LVT U3166 ( .A1(n3380), .A2(wdata[27]), .A3(n3379), .A4(
        \regs[27][27] ), .Y(n1694) );
  AO22X1_LVT U3167 ( .A1(n3384), .A2(n3503), .A3(n3383), .A4(\regs[27][26] ), 
        .Y(n1693) );
  AO22X1_LVT U3168 ( .A1(n3384), .A2(wdata[25]), .A3(n3383), .A4(
        \regs[27][25] ), .Y(n1692) );
  AO22X1_LVT U3170 ( .A1(n3382), .A2(n3493), .A3(n3381), .A4(\regs[27][24] ), 
        .Y(n1691) );
  AO22X1_LVT U3171 ( .A1(n3380), .A2(n3497), .A3(n3379), .A4(\regs[27][23] ), 
        .Y(n1690) );
  AO22X1_LVT U3172 ( .A1(n3380), .A2(n3494), .A3(n3379), .A4(\regs[27][22] ), 
        .Y(n1689) );
  AO22X1_LVT U3173 ( .A1(n3382), .A2(wdata[21]), .A3(n3381), .A4(
        \regs[27][21] ), .Y(n1688) );
  AO22X1_LVT U3174 ( .A1(n3380), .A2(n3483), .A3(n3379), .A4(\regs[27][20] ), 
        .Y(n1687) );
  AO22X1_LVT U3175 ( .A1(n3380), .A2(n3496), .A3(n3379), .A4(\regs[27][19] ), 
        .Y(n1686) );
  AO22X1_LVT U3176 ( .A1(n3380), .A2(n3491), .A3(n3379), .A4(\regs[27][18] ), 
        .Y(n1685) );
  AO22X1_LVT U3177 ( .A1(n3380), .A2(wdata[17]), .A3(n3379), .A4(
        \regs[27][17] ), .Y(n1684) );
  AO22X1_LVT U3179 ( .A1(n3380), .A2(wdata[16]), .A3(n3379), .A4(
        \regs[27][16] ), .Y(n1683) );
  AO22X1_LVT U3180 ( .A1(n3380), .A2(n3495), .A3(n3379), .A4(\regs[27][15] ), 
        .Y(n1682) );
  AO22X1_LVT U3181 ( .A1(n3380), .A2(n3498), .A3(n3379), .A4(\regs[27][14] ), 
        .Y(n1681) );
  AO22X1_LVT U3182 ( .A1(n3380), .A2(n3502), .A3(n3379), .A4(\regs[27][13] ), 
        .Y(n1680) );
  AO22X1_LVT U3183 ( .A1(n3380), .A2(wdata[12]), .A3(n3379), .A4(
        \regs[27][12] ), .Y(n1679) );
  AO22X1_LVT U3184 ( .A1(n3380), .A2(wdata[11]), .A3(n3379), .A4(
        \regs[27][11] ), .Y(n1678) );
  AO22X1_LVT U3185 ( .A1(n3380), .A2(n3499), .A3(n3379), .A4(\regs[27][10] ), 
        .Y(n1677) );
  AO22X1_LVT U3186 ( .A1(n3384), .A2(wdata[9]), .A3(n3383), .A4(\regs[27][9] ), 
        .Y(n1676) );
  AO22X1_LVT U3188 ( .A1(n3382), .A2(wdata[8]), .A3(n3381), .A4(\regs[27][8] ), 
        .Y(n1675) );
  AO22X1_LVT U3189 ( .A1(n3382), .A2(wdata[7]), .A3(n3381), .A4(\regs[27][7] ), 
        .Y(n1674) );
  AO22X1_LVT U3190 ( .A1(n3382), .A2(wdata[6]), .A3(n3381), .A4(\regs[27][6] ), 
        .Y(n1673) );
  AO22X1_LVT U3191 ( .A1(n3382), .A2(wdata[5]), .A3(n3381), .A4(\regs[27][5] ), 
        .Y(n1672) );
  AO22X1_LVT U3192 ( .A1(n3382), .A2(wdata[4]), .A3(n3381), .A4(\regs[27][4] ), 
        .Y(n1671) );
  AO22X1_LVT U3193 ( .A1(n3382), .A2(wdata[3]), .A3(n3381), .A4(\regs[27][3] ), 
        .Y(n1670) );
  AO22X1_LVT U3194 ( .A1(n3382), .A2(wdata[2]), .A3(n3381), .A4(\regs[27][2] ), 
        .Y(n1669) );
  AO22X1_LVT U3196 ( .A1(n3382), .A2(wdata[1]), .A3(n3381), .A4(\regs[27][1] ), 
        .Y(n1668) );
  AO22X1_LVT U3197 ( .A1(n3382), .A2(wdata[0]), .A3(n3381), .A4(\regs[27][0] ), 
        .Y(n1667) );
  NAND4X0_LVT U3198 ( .A1(n3470), .A2(n3254), .A3(n3192), .A4(n3191), .Y(n3193) );
  AO22X1_LVT U3203 ( .A1(n3300), .A2(n3486), .A3(n3299), .A4(\regs[28][31] ), 
        .Y(n1666) );
  AO22X1_LVT U3204 ( .A1(n3300), .A2(wdata[30]), .A3(n3299), .A4(
        \regs[28][30] ), .Y(n1665) );
  AO22X1_LVT U3205 ( .A1(n3300), .A2(n3501), .A3(n3299), .A4(\regs[28][29] ), 
        .Y(n1664) );
  AO22X1_LVT U3206 ( .A1(n3300), .A2(n3500), .A3(n3299), .A4(\regs[28][28] ), 
        .Y(n1663) );
  AO22X1_LVT U3207 ( .A1(n3300), .A2(wdata[27]), .A3(n3299), .A4(
        \regs[28][27] ), .Y(n1662) );
  AO22X1_LVT U3208 ( .A1(n3300), .A2(n3503), .A3(n3299), .A4(\regs[28][26] ), 
        .Y(n1661) );
  AO22X1_LVT U3209 ( .A1(n3300), .A2(wdata[25]), .A3(n3299), .A4(
        \regs[28][25] ), .Y(n1660) );
  AO22X1_LVT U3211 ( .A1(n3302), .A2(n3493), .A3(n3301), .A4(\regs[28][24] ), 
        .Y(n1659) );
  AO22X1_LVT U3212 ( .A1(n3302), .A2(n3497), .A3(n3301), .A4(\regs[28][23] ), 
        .Y(n1658) );
  AO22X1_LVT U3213 ( .A1(n3302), .A2(n3494), .A3(n3301), .A4(\regs[28][22] ), 
        .Y(n1657) );
  AO22X1_LVT U3214 ( .A1(n3302), .A2(wdata[21]), .A3(n3301), .A4(
        \regs[28][21] ), .Y(n1656) );
  AO22X1_LVT U3215 ( .A1(n3302), .A2(n3483), .A3(n3301), .A4(\regs[28][20] ), 
        .Y(n1655) );
  AO22X1_LVT U3216 ( .A1(n3302), .A2(n3496), .A3(n3301), .A4(\regs[28][19] ), 
        .Y(n1654) );
  AO22X1_LVT U3217 ( .A1(n3302), .A2(n3491), .A3(n3301), .A4(\regs[28][18] ), 
        .Y(n1653) );
  AO22X1_LVT U3218 ( .A1(n3302), .A2(wdata[17]), .A3(n3301), .A4(
        \regs[28][17] ), .Y(n1652) );
  AO22X1_LVT U3220 ( .A1(n3300), .A2(wdata[16]), .A3(n3299), .A4(
        \regs[28][16] ), .Y(n1651) );
  AO22X1_LVT U3221 ( .A1(n3300), .A2(n3495), .A3(n3299), .A4(\regs[28][15] ), 
        .Y(n1650) );
  AO22X1_LVT U3222 ( .A1(n3300), .A2(n3498), .A3(n3299), .A4(\regs[28][14] ), 
        .Y(n1649) );
  AO22X1_LVT U3223 ( .A1(n3300), .A2(n3502), .A3(n3299), .A4(\regs[28][13] ), 
        .Y(n1648) );
  AO22X1_LVT U3224 ( .A1(n3300), .A2(wdata[12]), .A3(n3299), .A4(
        \regs[28][12] ), .Y(n1647) );
  AO22X1_LVT U3225 ( .A1(n3300), .A2(wdata[11]), .A3(n3299), .A4(
        \regs[28][11] ), .Y(n1646) );
  AO22X1_LVT U3226 ( .A1(n3300), .A2(n3499), .A3(n3299), .A4(\regs[28][10] ), 
        .Y(n1645) );
  AO22X1_LVT U3227 ( .A1(n3300), .A2(wdata[9]), .A3(n3299), .A4(\regs[28][9] ), 
        .Y(n1644) );
  AO22X1_LVT U3229 ( .A1(n3300), .A2(wdata[8]), .A3(n3299), .A4(\regs[28][8] ), 
        .Y(n1643) );
  AO22X1_LVT U3230 ( .A1(n3300), .A2(wdata[7]), .A3(n3299), .A4(\regs[28][7] ), 
        .Y(n1642) );
  AO22X1_LVT U3231 ( .A1(n3300), .A2(wdata[6]), .A3(n3299), .A4(\regs[28][6] ), 
        .Y(n1641) );
  AO22X1_LVT U3232 ( .A1(n3300), .A2(wdata[5]), .A3(n3299), .A4(\regs[28][5] ), 
        .Y(n1640) );
  AO22X1_LVT U3233 ( .A1(n3300), .A2(wdata[4]), .A3(n3299), .A4(\regs[28][4] ), 
        .Y(n1639) );
  AO22X1_LVT U3234 ( .A1(n3302), .A2(wdata[3]), .A3(n3301), .A4(\regs[28][3] ), 
        .Y(n1638) );
  AO22X1_LVT U3235 ( .A1(n3302), .A2(wdata[2]), .A3(n3301), .A4(\regs[28][2] ), 
        .Y(n1637) );
  AO22X1_LVT U3237 ( .A1(n3302), .A2(wdata[1]), .A3(n3301), .A4(\regs[28][1] ), 
        .Y(n1636) );
  AO22X1_LVT U3238 ( .A1(n3302), .A2(wdata[0]), .A3(n3301), .A4(\regs[28][0] ), 
        .Y(n1635) );
  AO22X1_LVT U3244 ( .A1(n3324), .A2(n3486), .A3(n3323), .A4(\regs[29][31] ), 
        .Y(n1634) );
  AO22X1_LVT U3245 ( .A1(n3324), .A2(wdata[30]), .A3(n3323), .A4(
        \regs[29][30] ), .Y(n1633) );
  AO22X1_LVT U3246 ( .A1(n3324), .A2(n3501), .A3(n3323), .A4(\regs[29][29] ), 
        .Y(n1632) );
  AO22X1_LVT U3247 ( .A1(n3324), .A2(n3500), .A3(n3323), .A4(\regs[29][28] ), 
        .Y(n1631) );
  AO22X1_LVT U3248 ( .A1(n3324), .A2(wdata[27]), .A3(n3323), .A4(
        \regs[29][27] ), .Y(n1630) );
  AO22X1_LVT U3249 ( .A1(n3324), .A2(n3503), .A3(n3323), .A4(\regs[29][26] ), 
        .Y(n1629) );
  AO22X1_LVT U3250 ( .A1(n3324), .A2(wdata[25]), .A3(n3323), .A4(
        \regs[29][25] ), .Y(n1628) );
  AO22X1_LVT U3252 ( .A1(n3324), .A2(n3493), .A3(n3323), .A4(\regs[29][24] ), 
        .Y(n1627) );
  AO22X1_LVT U3253 ( .A1(n3324), .A2(n3497), .A3(n3323), .A4(\regs[29][23] ), 
        .Y(n1626) );
  AO22X1_LVT U3254 ( .A1(n3324), .A2(n3494), .A3(n3323), .A4(\regs[29][22] ), 
        .Y(n1625) );
  AO22X1_LVT U3255 ( .A1(n3328), .A2(wdata[21]), .A3(n3327), .A4(
        \regs[29][21] ), .Y(n1624) );
  AO22X1_LVT U3256 ( .A1(n3324), .A2(n3483), .A3(n3323), .A4(\regs[29][20] ), 
        .Y(n1623) );
  AO22X1_LVT U3257 ( .A1(n3324), .A2(n3496), .A3(n3323), .A4(\regs[29][19] ), 
        .Y(n1622) );
  AO22X1_LVT U3258 ( .A1(n3324), .A2(n3491), .A3(n3323), .A4(\regs[29][18] ), 
        .Y(n1621) );
  AO22X1_LVT U3259 ( .A1(n3328), .A2(wdata[17]), .A3(n3327), .A4(
        \regs[29][17] ), .Y(n1620) );
  AO22X1_LVT U3261 ( .A1(n3326), .A2(wdata[16]), .A3(n3325), .A4(
        \regs[29][16] ), .Y(n1619) );
  AO22X1_LVT U3262 ( .A1(n3326), .A2(n3495), .A3(n3325), .A4(\regs[29][15] ), 
        .Y(n1618) );
  AO22X1_LVT U3263 ( .A1(n3324), .A2(n3498), .A3(n3323), .A4(\regs[29][14] ), 
        .Y(n1617) );
  AO22X1_LVT U3264 ( .A1(n3326), .A2(n3502), .A3(n3325), .A4(\regs[29][13] ), 
        .Y(n1616) );
  AO22X1_LVT U3265 ( .A1(n3326), .A2(wdata[12]), .A3(n3325), .A4(
        \regs[29][12] ), .Y(n1615) );
  AO22X1_LVT U3266 ( .A1(n3324), .A2(wdata[11]), .A3(n3323), .A4(
        \regs[29][11] ), .Y(n1614) );
  AO22X1_LVT U3267 ( .A1(n3326), .A2(n3499), .A3(n3325), .A4(\regs[29][10] ), 
        .Y(n1613) );
  AO22X1_LVT U3268 ( .A1(n3324), .A2(wdata[9]), .A3(n3323), .A4(\regs[29][9] ), 
        .Y(n1612) );
  AO22X1_LVT U3270 ( .A1(n3328), .A2(wdata[8]), .A3(n3327), .A4(\regs[29][8] ), 
        .Y(n1611) );
  AO22X1_LVT U3271 ( .A1(n3328), .A2(wdata[7]), .A3(n3327), .A4(\regs[29][7] ), 
        .Y(n1610) );
  AO22X1_LVT U3272 ( .A1(n3328), .A2(wdata[6]), .A3(n3327), .A4(\regs[29][6] ), 
        .Y(n1609) );
  AO22X1_LVT U3273 ( .A1(n3328), .A2(wdata[5]), .A3(n3327), .A4(\regs[29][5] ), 
        .Y(n1608) );
  AO22X1_LVT U3274 ( .A1(n3328), .A2(wdata[4]), .A3(n3327), .A4(\regs[29][4] ), 
        .Y(n1607) );
  AO22X1_LVT U3275 ( .A1(n3328), .A2(wdata[3]), .A3(n3327), .A4(\regs[29][3] ), 
        .Y(n1606) );
  AO22X1_LVT U3276 ( .A1(n3328), .A2(wdata[2]), .A3(n3327), .A4(\regs[29][2] ), 
        .Y(n1605) );
  AO22X1_LVT U3278 ( .A1(n3328), .A2(wdata[1]), .A3(n3327), .A4(\regs[29][1] ), 
        .Y(n1604) );
  AO22X1_LVT U3279 ( .A1(n3328), .A2(wdata[0]), .A3(n3327), .A4(\regs[29][0] ), 
        .Y(n1603) );
  NAND3X0_LVT U3280 ( .A1(n3470), .A2(n3212), .A3(n3254), .Y(n3213) );
  AO22X1_LVT U3285 ( .A1(n3320), .A2(n3486), .A3(n3319), .A4(\regs[30][31] ), 
        .Y(n1602) );
  AO22X1_LVT U3286 ( .A1(n3322), .A2(wdata[30]), .A3(n3321), .A4(
        \regs[30][30] ), .Y(n1601) );
  AO22X1_LVT U3287 ( .A1(n3320), .A2(n3501), .A3(n3319), .A4(\regs[30][29] ), 
        .Y(n1600) );
  AO22X1_LVT U3288 ( .A1(n3322), .A2(n3500), .A3(n3321), .A4(\regs[30][28] ), 
        .Y(n1599) );
  AO22X1_LVT U3289 ( .A1(n3322), .A2(wdata[27]), .A3(n3321), .A4(
        \regs[30][27] ), .Y(n1598) );
  AO22X1_LVT U3290 ( .A1(n3320), .A2(n3503), .A3(n3319), .A4(\regs[30][26] ), 
        .Y(n1597) );
  AO22X1_LVT U3291 ( .A1(n3322), .A2(wdata[25]), .A3(n3321), .A4(
        \regs[30][25] ), .Y(n1596) );
  AO22X1_LVT U3293 ( .A1(n3320), .A2(n3493), .A3(n3319), .A4(\regs[30][24] ), 
        .Y(n1595) );
  AO22X1_LVT U3294 ( .A1(n3320), .A2(n3497), .A3(n3319), .A4(\regs[30][23] ), 
        .Y(n1594) );
  AO22X1_LVT U3295 ( .A1(n3320), .A2(n3494), .A3(n3319), .A4(\regs[30][22] ), 
        .Y(n1593) );
  AO22X1_LVT U3296 ( .A1(n3320), .A2(wdata[21]), .A3(n3319), .A4(
        \regs[30][21] ), .Y(n1592) );
  AO22X1_LVT U3297 ( .A1(n3322), .A2(n3483), .A3(n3321), .A4(\regs[30][20] ), 
        .Y(n1591) );
  AO22X1_LVT U3298 ( .A1(n3320), .A2(n3496), .A3(n3319), .A4(\regs[30][19] ), 
        .Y(n1590) );
  AO22X1_LVT U3299 ( .A1(n3320), .A2(n3491), .A3(n3319), .A4(\regs[30][18] ), 
        .Y(n1589) );
  AO22X1_LVT U3300 ( .A1(n3320), .A2(wdata[17]), .A3(n3319), .A4(
        \regs[30][17] ), .Y(n1588) );
  AO22X1_LVT U3302 ( .A1(n3322), .A2(wdata[16]), .A3(n3321), .A4(
        \regs[30][16] ), .Y(n1587) );
  AO22X1_LVT U3303 ( .A1(n3320), .A2(n3495), .A3(n3319), .A4(\regs[30][15] ), 
        .Y(n1586) );
  AO22X1_LVT U3304 ( .A1(n3322), .A2(n3498), .A3(n3321), .A4(\regs[30][14] ), 
        .Y(n1585) );
  AO22X1_LVT U3305 ( .A1(n3322), .A2(n3502), .A3(n3321), .A4(\regs[30][13] ), 
        .Y(n1584) );
  AO22X1_LVT U3306 ( .A1(n3320), .A2(wdata[12]), .A3(n3319), .A4(
        \regs[30][12] ), .Y(n1583) );
  AO22X1_LVT U3307 ( .A1(n3322), .A2(wdata[11]), .A3(n3321), .A4(
        \regs[30][11] ), .Y(n1582) );
  AO22X1_LVT U3308 ( .A1(n3320), .A2(n3499), .A3(n3319), .A4(\regs[30][10] ), 
        .Y(n1581) );
  AO22X1_LVT U3309 ( .A1(n3322), .A2(wdata[9]), .A3(n3321), .A4(\regs[30][9] ), 
        .Y(n1580) );
  AO22X1_LVT U3311 ( .A1(n3322), .A2(wdata[8]), .A3(n3321), .A4(\regs[30][8] ), 
        .Y(n1579) );
  AO22X1_LVT U3312 ( .A1(n3322), .A2(wdata[7]), .A3(n3321), .A4(\regs[30][7] ), 
        .Y(n1578) );
  AO22X1_LVT U3313 ( .A1(n3322), .A2(wdata[6]), .A3(n3321), .A4(\regs[30][6] ), 
        .Y(n1577) );
  AO22X1_LVT U3314 ( .A1(n3322), .A2(wdata[5]), .A3(n3321), .A4(\regs[30][5] ), 
        .Y(n1576) );
  AO22X1_LVT U3315 ( .A1(n3322), .A2(wdata[4]), .A3(n3321), .A4(\regs[30][4] ), 
        .Y(n1575) );
  AO22X1_LVT U3316 ( .A1(n3322), .A2(wdata[3]), .A3(n3321), .A4(\regs[30][3] ), 
        .Y(n1574) );
  AO22X1_LVT U3317 ( .A1(n3322), .A2(wdata[2]), .A3(n3321), .A4(\regs[30][2] ), 
        .Y(n1573) );
  AO22X1_LVT U3319 ( .A1(n3322), .A2(wdata[1]), .A3(n3321), .A4(\regs[30][1] ), 
        .Y(n1572) );
  AO22X1_LVT U3320 ( .A1(n3322), .A2(wdata[0]), .A3(n3321), .A4(\regs[30][0] ), 
        .Y(n1571) );
  NAND3X0_LVT U3321 ( .A1(n3470), .A2(n3255), .A3(n3254), .Y(n3256) );
  AO22X1_LVT U3326 ( .A1(n3304), .A2(n3486), .A3(n3303), .A4(\regs[31][31] ), 
        .Y(n1570) );
  AO22X1_LVT U3327 ( .A1(n3304), .A2(wdata[30]), .A3(n3303), .A4(
        \regs[31][30] ), .Y(n1569) );
  AO22X1_LVT U3328 ( .A1(n3304), .A2(n3501), .A3(n3303), .A4(\regs[31][29] ), 
        .Y(n1568) );
  AO22X1_LVT U3329 ( .A1(n3304), .A2(n3500), .A3(n3303), .A4(\regs[31][28] ), 
        .Y(n1567) );
  AO22X1_LVT U3330 ( .A1(n3304), .A2(wdata[27]), .A3(n3303), .A4(
        \regs[31][27] ), .Y(n1566) );
  AO22X1_LVT U3331 ( .A1(n3304), .A2(n3503), .A3(n3303), .A4(\regs[31][26] ), 
        .Y(n1565) );
  AO22X1_LVT U3332 ( .A1(n3304), .A2(wdata[25]), .A3(n3303), .A4(
        \regs[31][25] ), .Y(n1564) );
  AO22X1_LVT U3334 ( .A1(n3306), .A2(n3493), .A3(n3305), .A4(\regs[31][24] ), 
        .Y(n1563) );
  AO22X1_LVT U3335 ( .A1(n3306), .A2(n3497), .A3(n3305), .A4(\regs[31][23] ), 
        .Y(n1562) );
  AO22X1_LVT U3336 ( .A1(n3304), .A2(n3494), .A3(n3303), .A4(\regs[31][22] ), 
        .Y(n1561) );
  AO22X1_LVT U3337 ( .A1(n3306), .A2(wdata[21]), .A3(n3305), .A4(
        \regs[31][21] ), .Y(n1560) );
  AO22X1_LVT U3338 ( .A1(n3306), .A2(n3483), .A3(n3305), .A4(\regs[31][20] ), 
        .Y(n1559) );
  AO22X1_LVT U3339 ( .A1(n3306), .A2(n3496), .A3(n3305), .A4(\regs[31][19] ), 
        .Y(n1558) );
  AO22X1_LVT U3340 ( .A1(n3304), .A2(n3491), .A3(n3303), .A4(\regs[31][18] ), 
        .Y(n1557) );
  AO22X1_LVT U3341 ( .A1(n3304), .A2(wdata[17]), .A3(n3303), .A4(
        \regs[31][17] ), .Y(n1556) );
  AO22X1_LVT U3343 ( .A1(n3304), .A2(wdata[16]), .A3(n3303), .A4(
        \regs[31][16] ), .Y(n1555) );
  AO22X1_LVT U3344 ( .A1(n3304), .A2(n3495), .A3(n3303), .A4(\regs[31][15] ), 
        .Y(n1554) );
  AO22X1_LVT U3345 ( .A1(n3304), .A2(n3498), .A3(n3303), .A4(\regs[31][14] ), 
        .Y(n1553) );
  AO22X1_LVT U3346 ( .A1(n3304), .A2(n3502), .A3(n3303), .A4(\regs[31][13] ), 
        .Y(n1552) );
  AO22X1_LVT U3347 ( .A1(n3304), .A2(wdata[12]), .A3(n3303), .A4(
        \regs[31][12] ), .Y(n1551) );
  AO22X1_LVT U3348 ( .A1(n3304), .A2(wdata[11]), .A3(n3303), .A4(
        \regs[31][11] ), .Y(n1550) );
  AO22X1_LVT U3349 ( .A1(n3304), .A2(n3499), .A3(n3303), .A4(\regs[31][10] ), 
        .Y(n1549) );
  AO22X1_LVT U3350 ( .A1(n3304), .A2(wdata[9]), .A3(n3303), .A4(\regs[31][9] ), 
        .Y(n1548) );
  AO22X1_LVT U3352 ( .A1(n3306), .A2(wdata[8]), .A3(n3305), .A4(\regs[31][8] ), 
        .Y(n1547) );
  AO22X1_LVT U3353 ( .A1(n3306), .A2(wdata[7]), .A3(n3305), .A4(\regs[31][7] ), 
        .Y(n1546) );
  AO22X1_LVT U3354 ( .A1(n3306), .A2(wdata[6]), .A3(n3305), .A4(\regs[31][6] ), 
        .Y(n1545) );
  AO22X1_LVT U3355 ( .A1(n3306), .A2(wdata[5]), .A3(n3305), .A4(\regs[31][5] ), 
        .Y(n1544) );
  AO22X1_LVT U3356 ( .A1(n3306), .A2(wdata[4]), .A3(n3305), .A4(\regs[31][4] ), 
        .Y(n1543) );
  AO22X1_LVT U3357 ( .A1(n3306), .A2(wdata[3]), .A3(n3305), .A4(\regs[31][3] ), 
        .Y(n1542) );
  AO22X1_LVT U3358 ( .A1(n3306), .A2(wdata[2]), .A3(n3305), .A4(\regs[31][2] ), 
        .Y(n1541) );
  AO22X1_LVT U3360 ( .A1(n3306), .A2(wdata[1]), .A3(n3305), .A4(\regs[31][1] ), 
        .Y(n1540) );
  AO22X1_LVT U3361 ( .A1(n3306), .A2(wdata[0]), .A3(n3305), .A4(\regs[31][0] ), 
        .Y(n1539) );
  AND2X4_LVT U1041 ( .A1(n959), .A2(n962), .Y(n960) );
  AND2X4_LVT U152 ( .A1(n78), .A2(n77), .Y(n79) );
  AND2X4_LVT U1044 ( .A1(n962), .A2(n961), .Y(n963) );
  AND2X4_LVT U24 ( .A1(n77), .A2(n76), .Y(n8) );
  AND2X4_LVT U1147 ( .A1(n1013), .A2(n1019), .Y(n1014) );
  NAND2X2_LVT U2051 ( .A1(n3202), .A2(n2955), .Y(n2905) );
  NAND2X2_LVT U2093 ( .A1(n2955), .A2(n3212), .Y(n2914) );
  NAND2X4_LVT U2456 ( .A1(n3212), .A2(n3030), .Y(n3021) );
  NAND2X2_LVT U2497 ( .A1(n3255), .A2(n3030), .Y(n3031) );
  NAND2X0_LVT U2786 ( .A1(n3212), .A2(n3105), .Y(n3096) );
  NAND2X2_LVT U2827 ( .A1(n3255), .A2(n3105), .Y(n3106) );
  NAND3X2_LVT U2374 ( .A1(n3030), .A2(n3192), .A3(n3191), .Y(n3003) );
  NAND2X0_LVT U3157 ( .A1(n3255), .A2(n3181), .Y(n3182) );
  NAND3X0_LVT U2290 ( .A1(n3470), .A2(n2992), .A3(n3212), .Y(n2983) );
  NAND3X2_LVT U2620 ( .A1(n3470), .A2(n3212), .A3(n3067), .Y(n3058) );
  NAND3X0_LVT U2909 ( .A1(n3470), .A2(n3202), .A3(n3142), .Y(n3124) );
  NAND3X2_LVT U2991 ( .A1(n3470), .A2(n3255), .A3(n3142), .Y(n3143) );
  NAND3X2_LVT U3034 ( .A1(n3181), .A2(n3192), .A3(n3191), .Y(n3154) );
  NAND3X2_LVT U3239 ( .A1(n3470), .A2(n3202), .A3(n3254), .Y(n3203) );
  AND2X2_LVT U2134 ( .A1(waddr[1]), .A2(waddr[0]), .Y(n3255) );
  INVX2_LVT U2 ( .A(rst), .Y(n3297) );
  INVX1_LVT U4 ( .A(waddr[2]), .Y(n3298) );
  NBUFFX8_LVT U6 ( .A(n3193), .Y(n3299) );
  INVX4_LVT U15 ( .A(n3299), .Y(n3300) );
  NBUFFX4_LVT U25 ( .A(n3193), .Y(n3301) );
  INVX4_LVT U26 ( .A(n3301), .Y(n3302) );
  NBUFFX8_LVT U30 ( .A(n3256), .Y(n3303) );
  INVX4_LVT U31 ( .A(n3303), .Y(n3304) );
  NBUFFX4_LVT U35 ( .A(n3256), .Y(n3305) );
  INVX2_LVT U38 ( .A(n3305), .Y(n3306) );
  NBUFFX4_LVT U39 ( .A(n3115), .Y(n3307) );
  INVX2_LVT U43 ( .A(n3307), .Y(n3308) );
  INVX4_LVT U51 ( .A(n3309), .Y(n3310) );
  NBUFFX8_LVT U56 ( .A(n3040), .Y(n3311) );
  INVX4_LVT U60 ( .A(n3311), .Y(n3312) );
  NBUFFX4_LVT U61 ( .A(n3040), .Y(n3313) );
  INVX4_LVT U64 ( .A(n3313), .Y(n3314) );
  NBUFFX8_LVT U65 ( .A(n2965), .Y(n3315) );
  INVX4_LVT U68 ( .A(n3315), .Y(n3316) );
  NBUFFX4_LVT U69 ( .A(n2965), .Y(n3317) );
  INVX4_LVT U71 ( .A(n3317), .Y(n3318) );
  NBUFFX4_LVT U72 ( .A(n3213), .Y(n3319) );
  INVX2_LVT U75 ( .A(n3319), .Y(n3320) );
  NBUFFX4_LVT U76 ( .A(n3213), .Y(n3321) );
  INVX4_LVT U78 ( .A(n3321), .Y(n3322) );
  NBUFFX4_LVT U79 ( .A(n3203), .Y(n3323) );
  INVX2_LVT U82 ( .A(n3323), .Y(n3324) );
  NBUFFX4_LVT U83 ( .A(n3203), .Y(n3325) );
  INVX1_LVT U85 ( .A(n3325), .Y(n3326) );
  NBUFFX4_LVT U86 ( .A(n3203), .Y(n3327) );
  INVX2_LVT U91 ( .A(n3327), .Y(n3328) );
  NBUFFX4_LVT U92 ( .A(n3154), .Y(n3329) );
  INVX2_LVT U94 ( .A(n3329), .Y(n3330) );
  NBUFFX4_LVT U95 ( .A(n3154), .Y(n3331) );
  NBUFFX4_LVT U99 ( .A(n3143), .Y(n3333) );
  INVX2_LVT U101 ( .A(n3333), .Y(n3334) );
  NBUFFX4_LVT U102 ( .A(n3143), .Y(n3335) );
  INVX2_LVT U105 ( .A(n3335), .Y(n3336) );
  NBUFFX4_LVT U106 ( .A(n3143), .Y(n3337) );
  INVX1_LVT U108 ( .A(n3337), .Y(n3338) );
  NBUFFX4_LVT U109 ( .A(n3133), .Y(n3339) );
  INVX4_LVT U112 ( .A(n3339), .Y(n3340) );
  NBUFFX4_LVT U113 ( .A(n3133), .Y(n3341) );
  INVX4_LVT U115 ( .A(n3341), .Y(n3342) );
  NBUFFX4_LVT U116 ( .A(n3124), .Y(n3343) );
  INVX2_LVT U120 ( .A(n3343), .Y(n3344) );
  NBUFFX4_LVT U121 ( .A(n3124), .Y(n3345) );
  INVX2_LVT U123 ( .A(n3345), .Y(n3346) );
  INVX1_LVT U124 ( .A(n3348), .Y(n3347) );
  INVX2_LVT U131 ( .A(n3348), .Y(n3351) );
  NBUFFX4_LVT U134 ( .A(n3058), .Y(n3352) );
  INVX4_LVT U135 ( .A(n3352), .Y(n3353) );
  NBUFFX4_LVT U137 ( .A(n3058), .Y(n3354) );
  INVX1_LVT U138 ( .A(n3354), .Y(n3355) );
  NBUFFX4_LVT U141 ( .A(n3058), .Y(n3356) );
  INVX2_LVT U142 ( .A(n3356), .Y(n3357) );
  NBUFFX8_LVT U144 ( .A(n3049), .Y(n3358) );
  INVX4_LVT U145 ( .A(n3358), .Y(n3359) );
  NBUFFX4_LVT U150 ( .A(n3049), .Y(n3360) );
  INVX4_LVT U153 ( .A(n3360), .Y(n3361) );
  INVX1_LVT U154 ( .A(n3363), .Y(n3362) );
  INVX2_LVT U160 ( .A(n3363), .Y(n3364) );
  NBUFFX4_LVT U170 ( .A(n2983), .Y(n3367) );
  INVX2_LVT U173 ( .A(n3367), .Y(n3368) );
  NBUFFX4_LVT U175 ( .A(n2983), .Y(n3369) );
  INVX2_LVT U178 ( .A(n3369), .Y(n3370) );
  NBUFFX4_LVT U181 ( .A(n2983), .Y(n3371) );
  INVX4_LVT U184 ( .A(n3371), .Y(n3372) );
  NBUFFX4_LVT U190 ( .A(n2974), .Y(n3373) );
  INVX2_LVT U192 ( .A(n3373), .Y(n3374) );
  INVX2_LVT U195 ( .A(n3377), .Y(n3376) );
  NBUFFX4_LVT U198 ( .A(n3373), .Y(n3377) );
  INVX1_LVT U199 ( .A(n3377), .Y(n3378) );
  NBUFFX4_LVT U204 ( .A(n3182), .Y(n3379) );
  INVX4_LVT U205 ( .A(n3379), .Y(n3380) );
  NBUFFX4_LVT U207 ( .A(n3182), .Y(n3381) );
  INVX4_LVT U209 ( .A(n3381), .Y(n3382) );
  NBUFFX4_LVT U211 ( .A(n3182), .Y(n3383) );
  INVX1_LVT U214 ( .A(n3383), .Y(n3384) );
  NBUFFX4_LVT U216 ( .A(n3172), .Y(n3385) );
  INVX2_LVT U218 ( .A(n3385), .Y(n3386) );
  NBUFFX4_LVT U219 ( .A(n3172), .Y(n3387) );
  INVX2_LVT U223 ( .A(n3387), .Y(n3388) );
  NBUFFX4_LVT U225 ( .A(n3163), .Y(n3389) );
  INVX2_LVT U227 ( .A(n3389), .Y(n3390) );
  NBUFFX4_LVT U228 ( .A(n3163), .Y(n3391) );
  INVX4_LVT U230 ( .A(n3391), .Y(n3392) );
  NBUFFX4_LVT U231 ( .A(n3078), .Y(n3393) );
  INVX4_LVT U236 ( .A(n3393), .Y(n3394) );
  NBUFFX4_LVT U238 ( .A(n3078), .Y(n3395) );
  INVX2_LVT U240 ( .A(n3395), .Y(n3396) );
  NBUFFX4_LVT U243 ( .A(n3003), .Y(n3397) );
  INVX4_LVT U248 ( .A(n3397), .Y(n3398) );
  NBUFFX4_LVT U250 ( .A(n3003), .Y(n3399) );
  INVX1_LVT U253 ( .A(n3399), .Y(n3400) );
  NBUFFX4_LVT U258 ( .A(n3003), .Y(n3401) );
  INVX2_LVT U269 ( .A(n3401), .Y(n3402) );
  NBUFFX4_LVT U283 ( .A(n3106), .Y(n3403) );
  INVX2_LVT U284 ( .A(n3403), .Y(n3404) );
  NBUFFX4_LVT U286 ( .A(n3106), .Y(n3405) );
  INVX2_LVT U291 ( .A(n3405), .Y(n3406) );
  NBUFFX4_LVT U295 ( .A(n3106), .Y(n3407) );
  INVX2_LVT U300 ( .A(n3407), .Y(n3408) );
  INVX4_LVT U315 ( .A(n3409), .Y(n3410) );
  NBUFFX4_LVT U328 ( .A(n3096), .Y(n3411) );
  INVX4_LVT U354 ( .A(n3411), .Y(n3412) );
  NBUFFX4_LVT U375 ( .A(n3087), .Y(n3413) );
  INVX2_LVT U381 ( .A(n3413), .Y(n3414) );
  NBUFFX4_LVT U395 ( .A(n3087), .Y(n3415) );
  INVX2_LVT U399 ( .A(n3415), .Y(n3416) );
  NBUFFX4_LVT U409 ( .A(n3031), .Y(n3417) );
  NBUFFX4_LVT U440 ( .A(n3031), .Y(n3419) );
  INVX2_LVT U452 ( .A(n3419), .Y(n3420) );
  NBUFFX4_LVT U463 ( .A(n3031), .Y(n3421) );
  INVX1_LVT U499 ( .A(n3021), .Y(n3423) );
  NBUFFX4_LVT U516 ( .A(n3021), .Y(n3424) );
  NBUFFX4_LVT U543 ( .A(n3021), .Y(n3426) );
  INVX4_LVT U569 ( .A(n3426), .Y(n3427) );
  NBUFFX4_LVT U571 ( .A(n3012), .Y(n3428) );
  INVX2_LVT U596 ( .A(n3428), .Y(n3429) );
  NBUFFX4_LVT U597 ( .A(n3012), .Y(n3430) );
  INVX4_LVT U623 ( .A(n3430), .Y(n3431) );
  NBUFFX4_LVT U625 ( .A(n2956), .Y(n3432) );
  INVX4_LVT U650 ( .A(n3432), .Y(n3433) );
  NBUFFX4_LVT U676 ( .A(n2956), .Y(n3434) );
  INVX2_LVT U690 ( .A(n3434), .Y(n3435) );
  NBUFFX4_LVT U703 ( .A(n2914), .Y(n3436) );
  INVX2_LVT U729 ( .A(n3436), .Y(n3437) );
  NBUFFX4_LVT U755 ( .A(n2914), .Y(n3438) );
  INVX2_LVT U757 ( .A(n3438), .Y(n3439) );
  NBUFFX4_LVT U765 ( .A(n2914), .Y(n3440) );
  INVX1_LVT U783 ( .A(n3440), .Y(n3441) );
  NBUFFX4_LVT U800 ( .A(n2905), .Y(n3442) );
  INVX2_LVT U810 ( .A(n3442), .Y(n3443) );
  NBUFFX4_LVT U822 ( .A(n2905), .Y(n3444) );
  INVX2_LVT U837 ( .A(n3444), .Y(n3445) );
  NBUFFX4_LVT U863 ( .A(n2905), .Y(n3446) );
  INVX1_LVT U889 ( .A(n3446), .Y(n3447) );
  INVX1_LVT U915 ( .A(raddr2[3]), .Y(n3448) );
  INVX1_LVT U941 ( .A(raddr2[2]), .Y(n3449) );
  INVX1_LVT U967 ( .A(raddr1[2]), .Y(n3450) );
  INVX1_LVT U969 ( .A(raddr1[3]), .Y(n3451) );
  INVX1_LVT U994 ( .A(raddr1[4]), .Y(n3452) );
  AND2X4_LVT U114 ( .A1(n57), .A2(n55), .Y(n44) );
  AND2X4_LVT U107 ( .A1(n60), .A2(n41), .Y(n42) );
  AND2X4_LVT U111 ( .A1(n60), .A2(n55), .Y(n43) );
  AND2X4_LVT U63 ( .A1(n57), .A2(n59), .Y(n23) );
  AND2X4_LVT U90 ( .A1(n49), .A2(n53), .Y(n36) );
  AND2X4_LVT U77 ( .A1(n27), .A2(n49), .Y(n28) );
  AND2X4_LVT U100 ( .A1(n57), .A2(n53), .Y(n39) );
  AND2X4_LVT U97 ( .A1(n60), .A2(n62), .Y(n38) );
  AND2X4_LVT U136 ( .A1(n60), .A2(n59), .Y(n61) );
  AND2X4_LVT U67 ( .A1(n64), .A2(n41), .Y(n24) );
  AND2X4_LVT U119 ( .A1(n49), .A2(n59), .Y(n50) );
  AND2X4_LVT U29 ( .A1(n41), .A2(n57), .Y(n9) );
  AND2X4_LVT U37 ( .A1(n27), .A2(n57), .Y(n11) );
  AND2X4_LVT U34 ( .A1(n60), .A2(n27), .Y(n120) );
  AND2X4_LVT U126 ( .A1(n64), .A2(n53), .Y(n54) );
  AND2X4_LVT U140 ( .A1(n64), .A2(n62), .Y(n63) );
  AND2X4_LVT U50 ( .A1(n49), .A2(n62), .Y(n110) );
  AND2X4_LVT U104 ( .A1(n60), .A2(n53), .Y(n40) );
  AND2X4_LVT U47 ( .A1(n49), .A2(n55), .Y(n122) );
  AND2X4_LVT U74 ( .A1(n57), .A2(n62), .Y(n26) );
  AND2X4_LVT U42 ( .A1(n51), .A2(n49), .Y(n148) );
  AND2X4_LVT U84 ( .A1(n64), .A2(n59), .Y(n30) );
  AND2X4_LVT U129 ( .A1(n64), .A2(n55), .Y(n56) );
  AND2X4_LVT U122 ( .A1(n51), .A2(n64), .Y(n52) );
  AND2X4_LVT U93 ( .A1(n51), .A2(n57), .Y(n37) );
  AND2X4_LVT U55 ( .A1(n64), .A2(n27), .Y(n135) );
  AND2X4_LVT U70 ( .A1(n41), .A2(n49), .Y(n25) );
  AND2X4_LVT U1062 ( .A1(n1024), .A2(n1000), .Y(n969) );
  AND2X4_LVT U1151 ( .A1(n1026), .A2(n1023), .Y(n1015) );
  AND2X4_LVT U1059 ( .A1(n1026), .A2(n1000), .Y(n968) );
  AND2X4_LVT U1122 ( .A1(n1019), .A2(n1023), .Y(n997) );
  AND2X4_LVT U1110 ( .A1(n1024), .A2(n1016), .Y(n990) );
  AND2X4_LVT U1090 ( .A1(n1026), .A2(n1004), .Y(n982) );
  AND2X4_LVT U1161 ( .A1(n1026), .A2(n1021), .Y(n1022) );
  AND2X4_LVT U1129 ( .A1(n1011), .A2(n1000), .Y(n1001) );
  AND2X4_LVT U1115 ( .A1(n1019), .A2(n1016), .Y(n995) );
  AND2X4_LVT U1086 ( .A1(n1011), .A2(n1021), .Y(n981) );
  AND2X4_LVT U1054 ( .A1(n1024), .A2(n1021), .Y(n967) );
  AND2X4_LVT U1049 ( .A1(n1013), .A2(n1026), .Y(n965) );
  AND2X4_LVT U1144 ( .A1(n1011), .A2(n1018), .Y(n1012) );
  AND2X4_LVT U1165 ( .A1(n1024), .A2(n1023), .Y(n1025) );
  AND2X4_LVT U1158 ( .A1(n1019), .A2(n1018), .Y(n1020) );
  AND2X4_LVT U1132 ( .A1(n1019), .A2(n1004), .Y(n1002) );
  AND2X4_LVT U1154 ( .A1(n1026), .A2(n1016), .Y(n1017) );
  AND2X4_LVT U1082 ( .A1(n1024), .A2(n1004), .Y(n979) );
  AND2X4_LVT U1068 ( .A1(n1019), .A2(n1021), .Y(n972) );
  AND2X4_LVT U1136 ( .A1(n1011), .A2(n1016), .Y(n1003) );
  AND2X4_LVT U1106 ( .A1(n1024), .A2(n1018), .Y(n987) );
  AND2X4_LVT U1099 ( .A1(n1026), .A2(n1018), .Y(n985) );
  AND2X4_LVT U1118 ( .A1(n1019), .A2(n1000), .Y(n996) );
  AND2X4_LVT U1094 ( .A1(n1011), .A2(n1023), .Y(n983) );
  AND2X4_LVT U1139 ( .A1(n1011), .A2(n1004), .Y(n1005) );
  AND2X4_LVT U1125 ( .A1(n1013), .A2(n1024), .Y(n998) );
  AND4X4_LVT U143 ( .A1(raddr2[3]), .A2(raddr2[4]), .A3(raddr2[2]), .A4(n64), 
        .Y(n65) );
  AND4X4_LVT U133 ( .A1(raddr2[3]), .A2(raddr2[4]), .A3(raddr2[2]), .A4(n57), 
        .Y(n58) );
  AND4X4_LVT U59 ( .A1(raddr2[3]), .A2(raddr2[4]), .A3(raddr2[2]), .A4(n49), 
        .Y(n21) );
  AND4X4_LVT U81 ( .A1(raddr2[3]), .A2(raddr2[4]), .A3(raddr2[2]), .A4(n60), 
        .Y(n29) );
  DFFX2_LVT \regs_reg[17][30]  ( .D(n2017), .CLK(clk), .Q(\regs[17][30] ) );
  DFFX2_LVT \regs_reg[15][27]  ( .D(n2078), .CLK(clk), .Q(\regs[15][27] ) );
  DFFX2_LVT \regs_reg[24][30]  ( .D(n1793), .CLK(clk), .Q(\regs[24][30] ) );
  DFFX2_LVT \regs_reg[21][9]  ( .D(n1868), .CLK(clk), .Q(\regs[21][9] ) );
  DFFX2_LVT \regs_reg[21][30]  ( .D(n1889), .CLK(clk), .Q(\regs[21][30] ) );
  DFFX2_LVT \regs_reg[21][10]  ( .D(n1869), .CLK(clk), .Q(\regs[21][10] ) );
  DFFX2_LVT \regs_reg[26][9]  ( .D(n1708), .CLK(clk), .Q(\regs[26][9] ) );
  DFFX2_LVT \regs_reg[29][30]  ( .D(n1633), .CLK(clk), .Q(\regs[29][30] ) );
  DFFX2_LVT \regs_reg[2][23]  ( .D(n2490), .CLK(clk), .Q(\regs[2][23] ) );
  DFFX2_LVT \regs_reg[24][9]  ( .D(n1772), .CLK(clk), .Q(\regs[24][9] ) );
  DFFX2_LVT \regs_reg[24][10]  ( .D(n1773), .CLK(clk), .Q(\regs[24][10] ) );
  DFFX2_LVT \regs_reg[17][31]  ( .D(n2018), .CLK(clk), .Q(\regs[17][31] ) );
  DFFX2_LVT \regs_reg[31][11]  ( .D(n1550), .CLK(clk), .Q(\regs[31][11] ) );
  DFFX2_LVT \regs_reg[27][30]  ( .D(n1697), .CLK(clk), .Q(\regs[27][30] ) );
  DFFX2_LVT \regs_reg[2][19]  ( .D(n2486), .CLK(clk), .Q(\regs[2][19] ) );
  DFFX2_LVT \regs_reg[26][30]  ( .D(n1729), .CLK(clk), .Q(\regs[26][30] ) );
  DFFX2_LVT \regs_reg[26][10]  ( .D(n1709), .CLK(clk), .Q(\regs[26][10] ) );
  DFFX2_LVT \regs_reg[13][15]  ( .D(n2130), .CLK(clk), .Q(\regs[13][15] ) );
  DFFX2_LVT \regs_reg[24][26]  ( .D(n1789), .CLK(clk), .Q(\regs[24][26] ) );
  DFFX2_LVT \regs_reg[17][7]  ( .D(n1994), .CLK(clk), .Q(\regs[17][7] ) );
  DFFX2_LVT \regs_reg[26][16]  ( .D(n1715), .CLK(clk), .Q(\regs[26][16] ) );
  DFFX2_LVT \regs_reg[31][25]  ( .D(n1564), .CLK(clk), .Q(\regs[31][25] ) );
  DFFX2_LVT \regs_reg[26][31]  ( .D(n1730), .CLK(clk), .Q(\regs[26][31] ) );
  DFFX2_LVT \regs_reg[24][12]  ( .D(n1775), .CLK(clk), .Q(\regs[24][12] ) );
  DFFX2_LVT \regs_reg[2][24]  ( .D(n2491), .CLK(clk), .Q(\regs[2][24] ) );
  DFFX2_LVT \regs_reg[2][14]  ( .D(n2481), .CLK(clk), .Q(\regs[2][14] ) );
  DFFX2_LVT \regs_reg[17][10]  ( .D(n1997), .CLK(clk), .Q(\regs[17][10] ) );
  DFFX2_LVT \regs_reg[26][12]  ( .D(n1711), .CLK(clk), .Q(\regs[26][12] ) );
  DFFX2_LVT \regs_reg[13][14]  ( .D(n2129), .CLK(clk), .Q(\regs[13][14] ) );
  DFFX2_LVT \regs_reg[15][19]  ( .D(n2070), .CLK(clk), .Q(\regs[15][19] ) );
  DFFX2_LVT \regs_reg[21][12]  ( .D(n1871), .CLK(clk), .Q(\regs[21][12] ) );
  DFFX2_LVT \regs_reg[13][11]  ( .D(n2126), .CLK(clk), .Q(\regs[13][11] ) );
  DFFX2_LVT \regs_reg[26][5]  ( .D(n1704), .CLK(clk), .Q(\regs[26][5] ) );
  DFFX2_LVT \regs_reg[5][27]  ( .D(n2398), .CLK(clk), .Q(\regs[5][27] ) );
  DFFX2_LVT \regs_reg[24][31]  ( .D(n1794), .CLK(clk), .Q(\regs[24][31] ) );
  DFFX2_LVT \regs_reg[26][15]  ( .D(n1714), .CLK(clk), .Q(\regs[26][15] ) );
  DFFX2_LVT \regs_reg[26][17]  ( .D(n1716), .CLK(clk), .Q(\regs[26][17] ) );
  DFFX2_LVT \regs_reg[1][24]  ( .D(n2523), .CLK(clk), .Q(\regs[1][24] ) );
  DFFX2_LVT \regs_reg[31][29]  ( .D(n1568), .CLK(clk), .Q(\regs[31][29] ) );
  DFFX2_LVT \regs_reg[5][19]  ( .D(n2390), .CLK(clk), .Q(\regs[5][19] ) );
  DFFX2_LVT \regs_reg[21][28]  ( .D(n1887), .CLK(clk), .Q(\regs[21][28] ) );
  DFFX2_LVT \regs_reg[24][13]  ( .D(n1776), .CLK(clk), .Q(\regs[24][13] ) );
  DFFX2_LVT \regs_reg[28][17]  ( .D(n1652), .CLK(clk), .Q(\regs[28][17] ) );
  DFFX2_LVT \regs_reg[29][6]  ( .D(n1609), .CLK(clk), .Q(\regs[29][6] ) );
  DFFX2_LVT \regs_reg[24][28]  ( .D(n1791), .CLK(clk), .Q(\regs[24][28] ) );
  DFFX2_LVT \regs_reg[2][26]  ( .D(n2493), .CLK(clk), .Q(\regs[2][26] ) );
  DFFX2_LVT \regs_reg[21][29]  ( .D(n1888), .CLK(clk), .Q(\regs[21][29] ) );
  AND4X4_LVT U1168 ( .A1(raddr1[2]), .A2(raddr1[4]), .A3(raddr1[3]), .A4(n1026), .Y(n1027) );
  DFFX2_LVT \regs_reg[17][17]  ( .D(n2004), .CLK(clk), .Q(\regs[17][17] ) );
  DFFX2_LVT \regs_reg[21][4]  ( .D(n1863), .CLK(clk), .Q(\regs[21][4] ) );
  DFFX2_LVT \regs_reg[26][6]  ( .D(n1705), .CLK(clk), .Q(\regs[26][6] ) );
  DFFX2_LVT \regs_reg[2][27]  ( .D(n2494), .CLK(clk), .Q(\regs[2][27] ) );
  DFFX2_LVT \regs_reg[1][14]  ( .D(n2513), .CLK(clk), .Q(\regs[1][14] ) );
  DFFX2_LVT \regs_reg[21][6]  ( .D(n1865), .CLK(clk), .Q(\regs[21][6] ) );
  DFFX2_LVT \regs_reg[24][16]  ( .D(n1779), .CLK(clk), .Q(\regs[24][16] ) );
  DFFX2_LVT \regs_reg[1][18]  ( .D(n2517), .CLK(clk), .Q(\regs[1][18] ) );
  DFFX2_LVT \regs_reg[21][15]  ( .D(n1874), .CLK(clk), .Q(\regs[21][15] ) );
  DFFX2_LVT \regs_reg[7][28]  ( .D(n2335), .CLK(clk), .Q(\regs[7][28] ) );
  DFFX2_LVT \regs_reg[15][23]  ( .D(n2074), .CLK(clk), .Q(\regs[15][23] ) );
  DFFX2_LVT \regs_reg[29][9]  ( .D(n1612), .CLK(clk), .Q(\regs[29][9] ) );
  DFFX2_LVT \regs_reg[5][11]  ( .D(n2382), .CLK(clk), .Q(\regs[5][11] ) );
  DFFX2_LVT \regs_reg[1][5]  ( .D(n2504), .CLK(clk), .Q(\regs[1][5] ) );
  DFFX2_LVT \regs_reg[13][10]  ( .D(n2125), .CLK(clk), .Q(\regs[13][10] ) );
  DFFX2_LVT \regs_reg[15][14]  ( .D(n2065), .CLK(clk), .Q(\regs[15][14] ) );
  DFFX2_LVT \regs_reg[7][31]  ( .D(n2338), .CLK(clk), .Q(\regs[7][31] ) );
  DFFX2_LVT \regs_reg[13][12]  ( .D(n2127), .CLK(clk), .Q(\regs[13][12] ) );
  DFFX2_LVT \regs_reg[2][17]  ( .D(n2484), .CLK(clk), .Q(\regs[2][17] ) );
  DFFX2_LVT \regs_reg[24][29]  ( .D(n1792), .CLK(clk), .Q(\regs[24][29] ) );
  DFFX2_LVT \regs_reg[27][8]  ( .D(n1675), .CLK(clk), .Q(\regs[27][8] ) );
  DFFX2_LVT \regs_reg[10][26]  ( .D(n2237), .CLK(clk), .Q(\regs[10][26] ) );
  DFFX2_LVT \regs_reg[2][20]  ( .D(n2487), .CLK(clk), .Q(\regs[2][20] ) );
  DFFX2_LVT \regs_reg[23][29]  ( .D(n1824), .CLK(clk), .Q(\regs[23][29] ) );
  DFFX2_LVT \regs_reg[1][6]  ( .D(n2505), .CLK(clk), .Q(\regs[1][6] ) );
  DFFX2_LVT \regs_reg[17][19]  ( .D(n2006), .CLK(clk), .Q(\regs[17][19] ) );
  AND4X4_LVT U1076 ( .A1(raddr1[2]), .A2(raddr1[4]), .A3(raddr1[3]), .A4(n1019), .Y(n975) );
  DFFX2_LVT \regs_reg[17][6]  ( .D(n1993), .CLK(clk), .Q(\regs[17][6] ) );
  DFFX2_LVT \regs_reg[9][28]  ( .D(n2271), .CLK(clk), .Q(\regs[9][28] ) );
  DFFX2_LVT \regs_reg[5][24]  ( .D(n2395), .CLK(clk), .Q(\regs[5][24] ) );
  DFFX2_LVT \regs_reg[29][8]  ( .D(n1611), .CLK(clk), .Q(\regs[29][8] ) );
  DFFX2_LVT \regs_reg[2][25]  ( .D(n2492), .CLK(clk), .Q(\regs[2][25] ) );
  DFFX2_LVT \regs_reg[29][21]  ( .D(n1624), .CLK(clk), .Q(\regs[29][21] ) );
  DFFX2_LVT \regs_reg[1][26]  ( .D(n2525), .CLK(clk), .Q(\regs[1][26] ) );
  DFFX2_LVT \regs_reg[17][12]  ( .D(n1999), .CLK(clk), .Q(\regs[17][12] ) );
  AND4X4_LVT U1071 ( .A1(raddr1[2]), .A2(raddr1[4]), .A3(raddr1[3]), .A4(n1024), .Y(n973) );
  DFFX2_LVT \regs_reg[10][15]  ( .D(n2226), .CLK(clk), .Q(\regs[10][15] ) );
  DFFX2_LVT \regs_reg[5][20]  ( .D(n2391), .CLK(clk), .Q(\regs[5][20] ) );
  DFFX2_LVT \regs_reg[21][26]  ( .D(n1885), .CLK(clk), .Q(\regs[21][26] ) );
  DFFX2_LVT \regs_reg[17][13]  ( .D(n2000), .CLK(clk), .Q(\regs[17][13] ) );
  DFFX2_LVT \regs_reg[5][25]  ( .D(n2396), .CLK(clk), .Q(\regs[5][25] ) );
  DFFX2_LVT \regs_reg[7][19]  ( .D(n2326), .CLK(clk), .Q(\regs[7][19] ) );
  DFFX2_LVT \regs_reg[13][25]  ( .D(n2140), .CLK(clk), .Q(\regs[13][25] ) );
  DFFX2_LVT \regs_reg[24][15]  ( .D(n1778), .CLK(clk), .Q(\regs[24][15] ) );
  DFFX2_LVT \regs_reg[21][25]  ( .D(n1884), .CLK(clk), .Q(\regs[21][25] ) );
  DFFX2_LVT \regs_reg[26][4]  ( .D(n1703), .CLK(clk), .Q(\regs[26][4] ) );
  DFFX2_LVT \regs_reg[5][22]  ( .D(n2393), .CLK(clk), .Q(\regs[5][22] ) );
  DFFX2_LVT \regs_reg[21][7]  ( .D(n1866), .CLK(clk), .Q(\regs[21][7] ) );
  DFFX2_LVT \regs_reg[13][26]  ( .D(n2141), .CLK(clk), .Q(\regs[13][26] ) );
  DFFX2_LVT \regs_reg[21][31]  ( .D(n1890), .CLK(clk), .Q(\regs[21][31] ) );
  DFFX2_LVT \regs_reg[31][27]  ( .D(n1566), .CLK(clk), .Q(\regs[31][27] ) );
  DFFX2_LVT \regs_reg[26][7]  ( .D(n1706), .CLK(clk), .Q(\regs[26][7] ) );
  DFFX2_LVT \regs_reg[17][15]  ( .D(n2002), .CLK(clk), .Q(\regs[17][15] ) );
  DFFX2_LVT \regs_reg[2][18]  ( .D(n2485), .CLK(clk), .Q(\regs[2][18] ) );
  DFFX2_LVT \regs_reg[2][29]  ( .D(n2496), .CLK(clk), .Q(\regs[2][29] ) );
  DFFX2_LVT \regs_reg[13][16]  ( .D(n2131), .CLK(clk), .Q(\regs[13][16] ) );
  DFFX2_LVT \regs_reg[8][31]  ( .D(n2306), .CLK(clk), .Q(\regs[8][31] ) );
  DFFX2_LVT \regs_reg[8][28]  ( .D(n2303), .CLK(clk), .Q(\regs[8][28] ) );
  DFFX2_LVT \regs_reg[29][4]  ( .D(n1607), .CLK(clk), .Q(\regs[29][4] ) );
  DFFX2_LVT \regs_reg[30][9]  ( .D(n1580), .CLK(clk), .Q(\regs[30][9] ) );
  DFFX2_LVT \regs_reg[27][16]  ( .D(n1683), .CLK(clk), .Q(\regs[27][16] ) );
  DFFX2_LVT \regs_reg[29][28]  ( .D(n1631), .CLK(clk), .Q(\regs[29][28] ) );
  DFFX2_LVT \regs_reg[2][5]  ( .D(n2472), .CLK(clk), .Q(\regs[2][5] ) );
  DFFX2_LVT \regs_reg[2][21]  ( .D(n2488), .CLK(clk), .Q(\regs[2][21] ) );
  DFFX2_LVT \regs_reg[14][28]  ( .D(n2111), .CLK(clk), .Q(\regs[14][28] ) );
  DFFX2_LVT \regs_reg[21][13]  ( .D(n1872), .CLK(clk), .Q(\regs[21][13] ) );
  DFFX2_LVT \regs_reg[26][11]  ( .D(n1710), .CLK(clk), .Q(\regs[26][11] ) );
  DFFX2_LVT \regs_reg[21][5]  ( .D(n1864), .CLK(clk), .Q(\regs[21][5] ) );
  DFFX2_LVT \regs_reg[14][30]  ( .D(n2113), .CLK(clk), .Q(\regs[14][30] ) );
  DFFX2_LVT \regs_reg[15][24]  ( .D(n2075), .CLK(clk), .Q(\regs[15][24] ) );
  DFFX2_LVT \regs_reg[2][9]  ( .D(n2476), .CLK(clk), .Q(\regs[2][9] ) );
  DFFX2_LVT \regs_reg[29][5]  ( .D(n1608), .CLK(clk), .Q(\regs[29][5] ) );
  DFFX2_LVT \regs_reg[21][16]  ( .D(n1875), .CLK(clk), .Q(\regs[21][16] ) );
  DFFX2_LVT \regs_reg[27][6]  ( .D(n1673), .CLK(clk), .Q(\regs[27][6] ) );
  DFFX2_LVT \regs_reg[30][16]  ( .D(n1587), .CLK(clk), .Q(\regs[30][16] ) );
  DFFX2_LVT \regs_reg[10][14]  ( .D(n2225), .CLK(clk), .Q(\regs[10][14] ) );
  DFFX2_LVT \regs_reg[1][31]  ( .D(n2530), .CLK(clk), .Q(\regs[1][31] ) );
  DFFX2_LVT \regs_reg[30][7]  ( .D(n1578), .CLK(clk), .Q(\regs[30][7] ) );
  DFFX2_LVT \regs_reg[17][16]  ( .D(n2003), .CLK(clk), .Q(\regs[17][16] ) );
  DFFX2_LVT \regs_reg[1][20]  ( .D(n2519), .CLK(clk), .Q(\regs[1][20] ) );
  DFFX2_LVT \regs_reg[5][14]  ( .D(n2385), .CLK(clk), .Q(\regs[5][14] ) );
  DFFX2_LVT \regs_reg[15][9]  ( .D(n2060), .CLK(clk), .Q(\regs[15][9] ) );
  DFFX2_LVT \regs_reg[23][23]  ( .D(n1818), .CLK(clk), .Q(\regs[23][23] ) );
  DFFX2_LVT \regs_reg[24][14]  ( .D(n1777), .CLK(clk), .Q(\regs[24][14] ) );
  DFFX2_LVT \regs_reg[9][31]  ( .D(n2274), .CLK(clk), .Q(\regs[9][31] ) );
  DFFX2_LVT \regs_reg[15][11]  ( .D(n2062), .CLK(clk), .Q(\regs[15][11] ) );
  DFFX2_LVT \regs_reg[27][19]  ( .D(n1686), .CLK(clk), .Q(\regs[27][19] ) );
  DFFX2_LVT \regs_reg[17][8]  ( .D(n1995), .CLK(clk), .Q(\regs[17][8] ) );
  DFFX2_LVT \regs_reg[6][28]  ( .D(n2367), .CLK(clk), .Q(\regs[6][28] ) );
  DFFX2_LVT \regs_reg[15][25]  ( .D(n2076), .CLK(clk), .Q(\regs[15][25] ) );
  AND4X4_LVT U1102 ( .A1(raddr1[2]), .A2(raddr1[4]), .A3(raddr1[3]), .A4(n1011), .Y(n986) );
  DFFX2_LVT \regs_reg[15][20]  ( .D(n2071), .CLK(clk), .Q(\regs[15][20] ) );
  DFFX2_LVT \regs_reg[17][5]  ( .D(n1992), .CLK(clk), .Q(\regs[17][5] ) );
  DFFX2_LVT \regs_reg[2][15]  ( .D(n2482), .CLK(clk), .Q(\regs[2][15] ) );
  DFFX2_LVT \regs_reg[14][26]  ( .D(n2109), .CLK(clk), .Q(\regs[14][26] ) );
  DFFX2_LVT \regs_reg[26][29]  ( .D(n1728), .CLK(clk), .Q(\regs[26][29] ) );
  DFFX2_LVT \regs_reg[21][27]  ( .D(n1886), .CLK(clk), .Q(\regs[21][27] ) );
  DFFX2_LVT \regs_reg[27][15]  ( .D(n1682), .CLK(clk), .Q(\regs[27][15] ) );
  DFFX2_LVT \regs_reg[24][7]  ( .D(n1770), .CLK(clk), .Q(\regs[24][7] ) );
  DFFX2_LVT \regs_reg[14][31]  ( .D(n2114), .CLK(clk), .Q(\regs[14][31] ) );
  DFFX2_LVT \regs_reg[17][26]  ( .D(n2013), .CLK(clk), .Q(\regs[17][26] ) );
  DFFX2_LVT \regs_reg[15][26]  ( .D(n2077), .CLK(clk), .Q(\regs[15][26] ) );
  DFFX2_LVT \regs_reg[10][28]  ( .D(n2239), .CLK(clk), .Q(\regs[10][28] ) );
  DFFX2_LVT \regs_reg[23][17]  ( .D(n1812), .CLK(clk), .Q(\regs[23][17] ) );
  DFFX2_LVT \regs_reg[13][31]  ( .D(n2146), .CLK(clk), .Q(\regs[13][31] ) );
  DFFX2_LVT \regs_reg[1][23]  ( .D(n2522), .CLK(clk), .Q(\regs[1][23] ) );
  DFFX2_LVT \regs_reg[14][27]  ( .D(n2110), .CLK(clk), .Q(\regs[14][27] ) );
  DFFX2_LVT \regs_reg[24][5]  ( .D(n1768), .CLK(clk), .Q(\regs[24][5] ) );
  DFFX2_LVT \regs_reg[10][30]  ( .D(n2241), .CLK(clk), .Q(\regs[10][30] ) );
  DFFX2_LVT \regs_reg[30][4]  ( .D(n1575), .CLK(clk), .Q(\regs[30][4] ) );
  DFFX2_LVT \regs_reg[17][24]  ( .D(n2011), .CLK(clk), .Q(\regs[17][24] ) );
  DFFX2_LVT \regs_reg[31][26]  ( .D(n1565), .CLK(clk), .Q(\regs[31][26] ) );
  DFFX2_LVT \regs_reg[28][14]  ( .D(n1649), .CLK(clk), .Q(\regs[28][14] ) );
  DFFX2_LVT \regs_reg[17][9]  ( .D(n1996), .CLK(clk), .Q(\regs[17][9] ) );
  DFFX2_LVT \regs_reg[27][12]  ( .D(n1679), .CLK(clk), .Q(\regs[27][12] ) );
  DFFX2_LVT \regs_reg[31][15]  ( .D(n1554), .CLK(clk), .Q(\regs[31][15] ) );
  DFFX2_LVT \regs_reg[22][4]  ( .D(n1831), .CLK(clk), .Q(\regs[22][4] ) );
  DFFX2_LVT \regs_reg[2][28]  ( .D(n2495), .CLK(clk), .Q(\regs[2][28] ) );
  DFFX2_LVT \regs_reg[26][21]  ( .D(n1720), .CLK(clk), .Q(\regs[26][21] ) );
  DFFX2_LVT \regs_reg[7][29]  ( .D(n2336), .CLK(clk), .Q(\regs[7][29] ) );
  DFFX2_LVT \regs_reg[7][20]  ( .D(n2327), .CLK(clk), .Q(\regs[7][20] ) );
  DFFX2_LVT \regs_reg[26][8]  ( .D(n1707), .CLK(clk), .Q(\regs[26][8] ) );
  DFFX2_LVT \regs_reg[1][15]  ( .D(n2514), .CLK(clk), .Q(\regs[1][15] ) );
  DFFX2_LVT \regs_reg[22][6]  ( .D(n1833), .CLK(clk), .Q(\regs[22][6] ) );
  DFFX2_LVT \regs_reg[14][7]  ( .D(n2090), .CLK(clk), .Q(\regs[14][7] ) );
  DFFX2_LVT \regs_reg[29][7]  ( .D(n1610), .CLK(clk), .Q(\regs[29][7] ) );
  DFFX2_LVT \regs_reg[1][25]  ( .D(n2524), .CLK(clk), .Q(\regs[1][25] ) );
  DFFX2_LVT \regs_reg[15][29]  ( .D(n2080), .CLK(clk), .Q(\regs[15][29] ) );
  DFFX2_LVT \regs_reg[21][11]  ( .D(n1870), .CLK(clk), .Q(\regs[21][11] ) );
  DFFX2_LVT \regs_reg[6][17]  ( .D(n2356), .CLK(clk), .Q(\regs[6][17] ) );
  DFFX2_LVT \regs_reg[5][15]  ( .D(n2386), .CLK(clk), .Q(\regs[5][15] ) );
  DFFX2_LVT \regs_reg[13][30]  ( .D(n2145), .CLK(clk), .Q(\regs[13][30] ) );
  DFFX2_LVT \regs_reg[24][21]  ( .D(n1784), .CLK(clk), .Q(\regs[24][21] ) );
  DFFX2_LVT \regs_reg[27][29]  ( .D(n1696), .CLK(clk), .Q(\regs[27][29] ) );
  DFFX2_LVT \regs_reg[9][7]  ( .D(n2250), .CLK(clk), .Q(\regs[9][7] ) );
  DFFX2_LVT \regs_reg[7][23]  ( .D(n2330), .CLK(clk), .Q(\regs[7][23] ) );
  DFFX2_LVT \regs_reg[26][13]  ( .D(n1712), .CLK(clk), .Q(\regs[26][13] ) );
  DFFX2_LVT \regs_reg[19][14]  ( .D(n1937), .CLK(clk), .Q(\regs[19][14] ) );
  DFFX2_LVT \regs_reg[27][13]  ( .D(n1680), .CLK(clk), .Q(\regs[27][13] ) );
  DFFX2_LVT \regs_reg[1][9]  ( .D(n2508), .CLK(clk), .Q(\regs[1][9] ) );
  DFFX2_LVT \regs_reg[17][21]  ( .D(n2008), .CLK(clk), .Q(\regs[17][21] ) );
  DFFX2_LVT \regs_reg[15][12]  ( .D(n2063), .CLK(clk), .Q(\regs[15][12] ) );
  DFFX2_LVT \regs_reg[26][26]  ( .D(n1725), .CLK(clk), .Q(\regs[26][26] ) );
  DFFX2_LVT \regs_reg[21][14]  ( .D(n1873), .CLK(clk), .Q(\regs[21][14] ) );
  DFFX2_LVT \regs_reg[5][28]  ( .D(n2399), .CLK(clk), .Q(\regs[5][28] ) );
  DFFX2_LVT \regs_reg[7][25]  ( .D(n2332), .CLK(clk), .Q(\regs[7][25] ) );
  DFFX2_LVT \regs_reg[28][21]  ( .D(n1656), .CLK(clk), .Q(\regs[28][21] ) );
  DFFX2_LVT \regs_reg[15][8]  ( .D(n2059), .CLK(clk), .Q(\regs[15][8] ) );
  DFFX2_LVT \regs_reg[17][14]  ( .D(n2001), .CLK(clk), .Q(\regs[17][14] ) );
  DFFX2_LVT \regs_reg[24][11]  ( .D(n1774), .CLK(clk), .Q(\regs[24][11] ) );
  DFFX2_LVT \regs_reg[29][17]  ( .D(n1620), .CLK(clk), .Q(\regs[29][17] ) );
  DFFX2_LVT \regs_reg[26][25]  ( .D(n1724), .CLK(clk), .Q(\regs[26][25] ) );
  DFFX2_LVT \regs_reg[22][15]  ( .D(n1842), .CLK(clk), .Q(\regs[22][15] ) );
  DFFX2_LVT \regs_reg[15][31]  ( .D(n2082), .CLK(clk), .Q(\regs[15][31] ) );
  DFFX2_LVT \regs_reg[5][10]  ( .D(n2381), .CLK(clk), .Q(\regs[5][10] ) );
  DFFX2_LVT \regs_reg[29][27]  ( .D(n1630), .CLK(clk), .Q(\regs[29][27] ) );
  DFFX2_LVT \regs_reg[6][23]  ( .D(n2362), .CLK(clk), .Q(\regs[6][23] ) );
  DFFX2_LVT \regs_reg[30][29]  ( .D(n1600), .CLK(clk), .Q(\regs[30][29] ) );
  DFFX2_LVT \regs_reg[22][14]  ( .D(n1841), .CLK(clk), .Q(\regs[22][14] ) );
  DFFX2_LVT \regs_reg[9][5]  ( .D(n2248), .CLK(clk), .Q(\regs[9][5] ) );
  DFFX2_LVT \regs_reg[2][8]  ( .D(n2475), .CLK(clk), .Q(\regs[2][8] ) );
  DFFX2_LVT \regs_reg[29][25]  ( .D(n1628), .CLK(clk), .Q(\regs[29][25] ) );
  DFFX2_LVT \regs_reg[2][10]  ( .D(n2477), .CLK(clk), .Q(\regs[2][10] ) );
  DFFX2_LVT \regs_reg[10][25]  ( .D(n2236), .CLK(clk), .Q(\regs[10][25] ) );
  DFFX2_LVT \regs_reg[4][5]  ( .D(n2408), .CLK(clk), .Q(\regs[4][5] ) );
  DFFX2_LVT \regs_reg[17][25]  ( .D(n2012), .CLK(clk), .Q(\regs[17][25] ) );
  DFFX2_LVT \regs_reg[31][5]  ( .D(n1544), .CLK(clk), .Q(\regs[31][5] ) );
  DFFX2_LVT \regs_reg[31][10]  ( .D(n1549), .CLK(clk), .Q(\regs[31][10] ) );
  DFFX2_LVT \regs_reg[24][27]  ( .D(n1790), .CLK(clk), .Q(\regs[24][27] ) );
  DFFX2_LVT \regs_reg[28][4]  ( .D(n1639), .CLK(clk), .Q(\regs[28][4] ) );
  DFFX2_LVT \regs_reg[9][6]  ( .D(n2249), .CLK(clk), .Q(\regs[9][6] ) );
  DFFX2_LVT \regs_reg[3][25]  ( .D(n2460), .CLK(clk), .Q(\regs[3][25] ) );
  DFFX2_LVT \regs_reg[31][13]  ( .D(n1552), .CLK(clk), .Q(\regs[31][13] ) );
  DFFX2_LVT \regs_reg[8][27]  ( .D(n2302), .CLK(clk), .Q(\regs[8][27] ) );
  DFFX2_LVT \regs_reg[26][28]  ( .D(n1727), .CLK(clk), .Q(\regs[26][28] ) );
  DFFX2_LVT \regs_reg[2][16]  ( .D(n2483), .CLK(clk), .Q(\regs[2][16] ) );
  DFFX2_LVT \regs_reg[31][28]  ( .D(n1567), .CLK(clk), .Q(\regs[31][28] ) );
  DFFX2_LVT \regs_reg[9][15]  ( .D(n2258), .CLK(clk), .Q(\regs[9][15] ) );
  DFFX2_LVT \regs_reg[27][10]  ( .D(n1677), .CLK(clk), .Q(\regs[27][10] ) );
  DFFX2_LVT \regs_reg[30][13]  ( .D(n1584), .CLK(clk), .Q(\regs[30][13] ) );
  DFFX2_LVT \regs_reg[28][9]  ( .D(n1644), .CLK(clk), .Q(\regs[28][9] ) );
  DFFX2_LVT \regs_reg[27][11]  ( .D(n1678), .CLK(clk), .Q(\regs[27][11] ) );
  DFFX2_LVT \regs_reg[9][13]  ( .D(n2256), .CLK(clk), .Q(\regs[9][13] ) );
  DFFX2_LVT \regs_reg[17][22]  ( .D(n2009), .CLK(clk), .Q(\regs[17][22] ) );
  DFFX2_LVT \regs_reg[6][30]  ( .D(n2369), .CLK(clk), .Q(\regs[6][30] ) );
  DFFX2_LVT \regs_reg[22][17]  ( .D(n1844), .CLK(clk), .Q(\regs[22][17] ) );
  DFFX2_LVT \regs_reg[9][18]  ( .D(n2261), .CLK(clk), .Q(\regs[9][18] ) );
  DFFX2_LVT \regs_reg[10][23]  ( .D(n2234), .CLK(clk), .Q(\regs[10][23] ) );
  DFFX2_LVT \regs_reg[15][13]  ( .D(n2064), .CLK(clk), .Q(\regs[15][13] ) );
  DFFX2_LVT \regs_reg[29][3]  ( .D(n1606), .CLK(clk), .Q(\regs[29][3] ) );
  DFFX2_LVT \regs_reg[5][8]  ( .D(n2379), .CLK(clk), .Q(\regs[5][8] ) );
  DFFX2_LVT \regs_reg[21][8]  ( .D(n1867), .CLK(clk), .Q(\regs[21][8] ) );
  DFFX2_LVT \regs_reg[1][16]  ( .D(n2515), .CLK(clk), .Q(\regs[1][16] ) );
  DFFX2_LVT \regs_reg[2][11]  ( .D(n2478), .CLK(clk), .Q(\regs[2][11] ) );
  DFFX2_LVT \regs_reg[25][31]  ( .D(n1762), .CLK(clk), .Q(\regs[25][31] ) );
  DFFX2_LVT \regs_reg[10][11]  ( .D(n2222), .CLK(clk), .Q(\regs[10][11] ) );
  DFFX2_LVT \regs_reg[12][29]  ( .D(n2176), .CLK(clk), .Q(\regs[12][29] ) );
  DFFX2_LVT \regs_reg[5][31]  ( .D(n2402), .CLK(clk), .Q(\regs[5][31] ) );
  DFFX2_LVT \regs_reg[24][25]  ( .D(n1788), .CLK(clk), .Q(\regs[24][25] ) );
  DFFX2_LVT \regs_reg[10][20]  ( .D(n2231), .CLK(clk), .Q(\regs[10][20] ) );
  DFFX2_LVT \regs_reg[5][9]  ( .D(n2380), .CLK(clk), .Q(\regs[5][9] ) );
  DFFX2_LVT \regs_reg[31][14]  ( .D(n1553), .CLK(clk), .Q(\regs[31][14] ) );
  DFFX2_LVT \regs_reg[29][26]  ( .D(n1629), .CLK(clk), .Q(\regs[29][26] ) );
  DFFX2_LVT \regs_reg[30][22]  ( .D(n1593), .CLK(clk), .Q(\regs[30][22] ) );
  DFFX2_LVT \regs_reg[23][21]  ( .D(n1816), .CLK(clk), .Q(\regs[23][21] ) );
  DFFX2_LVT \regs_reg[13][5]  ( .D(n2120), .CLK(clk), .Q(\regs[13][5] ) );
  DFFX2_LVT \regs_reg[13][23]  ( .D(n2138), .CLK(clk), .Q(\regs[13][23] ) );
  DFFX2_LVT \regs_reg[2][31]  ( .D(n2498), .CLK(clk), .Q(\regs[2][31] ) );
  DFFX2_LVT \regs_reg[28][25]  ( .D(n1660), .CLK(clk), .Q(\regs[28][25] ) );
  DFFX2_LVT \regs_reg[31][31]  ( .D(n1570), .CLK(clk), .Q(\regs[31][31] ) );
  DFFX2_LVT \regs_reg[1][11]  ( .D(n2510), .CLK(clk), .Q(\regs[1][11] ) );
  DFFX2_LVT \regs_reg[15][30]  ( .D(n2081), .CLK(clk), .Q(\regs[15][30] ) );
  DFFX2_LVT \regs_reg[8][9]  ( .D(n2284), .CLK(clk), .Q(\regs[8][9] ) );
  DFFX2_LVT \regs_reg[1][8]  ( .D(n2507), .CLK(clk), .Q(\regs[1][8] ) );
  DFFX2_LVT \regs_reg[17][11]  ( .D(n1998), .CLK(clk), .Q(\regs[17][11] ) );
  DFFX2_LVT \regs_reg[5][30]  ( .D(n2401), .CLK(clk), .Q(\regs[5][30] ) );
  DFFX2_LVT \regs_reg[31][30]  ( .D(n1569), .CLK(clk), .Q(\regs[31][30] ) );
  DFFX2_LVT \regs_reg[23][27]  ( .D(n1822), .CLK(clk), .Q(\regs[23][27] ) );
  DFFX2_LVT \regs_reg[31][6]  ( .D(n1545), .CLK(clk), .Q(\regs[31][6] ) );
  DFFX2_LVT \regs_reg[2][30]  ( .D(n2497), .CLK(clk), .Q(\regs[2][30] ) );
  DFFX2_LVT \regs_reg[28][11]  ( .D(n1646), .CLK(clk), .Q(\regs[28][11] ) );
  DFFX2_LVT \regs_reg[2][6]  ( .D(n2473), .CLK(clk), .Q(\regs[2][6] ) );
  DFFX2_LVT \regs_reg[19][11]  ( .D(n1934), .CLK(clk), .Q(\regs[19][11] ) );
  DFFX2_LVT \regs_reg[20][21]  ( .D(n1912), .CLK(clk), .Q(\regs[20][21] ) );
  DFFX2_LVT \regs_reg[24][6]  ( .D(n1769), .CLK(clk), .Q(\regs[24][6] ) );
  DFFX2_LVT \regs_reg[7][30]  ( .D(n2337), .CLK(clk), .Q(\regs[7][30] ) );
  DFFX2_LVT \regs_reg[24][8]  ( .D(n1771), .CLK(clk), .Q(\regs[24][8] ) );
  DFFX2_LVT \regs_reg[14][11]  ( .D(n2094), .CLK(clk), .Q(\regs[14][11] ) );
  DFFX2_LVT \regs_reg[31][9]  ( .D(n1548), .CLK(clk), .Q(\regs[31][9] ) );
  DFFX2_LVT \regs_reg[14][4]  ( .D(n2087), .CLK(clk), .Q(\regs[14][4] ) );
  DFFX2_LVT \regs_reg[14][6]  ( .D(n2089), .CLK(clk), .Q(\regs[14][6] ) );
  DFFX2_LVT \regs_reg[25][25]  ( .D(n1756), .CLK(clk), .Q(\regs[25][25] ) );
  DFFX2_LVT \regs_reg[30][11]  ( .D(n1582), .CLK(clk), .Q(\regs[30][11] ) );
  DFFX2_LVT \regs_reg[16][7]  ( .D(n2026), .CLK(clk), .Q(\regs[16][7] ) );
  DFFX2_LVT \regs_reg[10][16]  ( .D(n2227), .CLK(clk), .Q(\regs[10][16] ) );
  DFFX2_LVT \regs_reg[7][21]  ( .D(n2328), .CLK(clk), .Q(\regs[7][21] ) );
  DFFX2_LVT \regs_reg[31][21]  ( .D(n1560), .CLK(clk), .Q(\regs[31][21] ) );
  DFFX2_LVT \regs_reg[15][15]  ( .D(n2066), .CLK(clk), .Q(\regs[15][15] ) );
  DFFX2_LVT \regs_reg[3][11]  ( .D(n2446), .CLK(clk), .Q(\regs[3][11] ) );
  DFFX2_LVT \regs_reg[18][25]  ( .D(n1980), .CLK(clk), .Q(\regs[18][25] ) );
  DFFX2_LVT \regs_reg[3][9]  ( .D(n2444), .CLK(clk), .Q(\regs[3][9] ) );
  DFFX2_LVT \regs_reg[5][12]  ( .D(n2383), .CLK(clk), .Q(\regs[5][12] ) );
  DFFX2_LVT \regs_reg[30][5]  ( .D(n1576), .CLK(clk), .Q(\regs[30][5] ) );
  DFFX2_LVT \regs_reg[5][3]  ( .D(n2374), .CLK(clk), .Q(\regs[5][3] ) );
  DFFX2_LVT \regs_reg[31][12]  ( .D(n1551), .CLK(clk), .Q(\regs[31][12] ) );
  DFFX2_LVT \regs_reg[9][9]  ( .D(n2252), .CLK(clk), .Q(\regs[9][9] ) );
  DFFX2_LVT \regs_reg[14][3]  ( .D(n2086), .CLK(clk), .Q(\regs[14][3] ) );
  DFFX2_LVT \regs_reg[9][11]  ( .D(n2254), .CLK(clk), .Q(\regs[9][11] ) );
  DFFX2_LVT \regs_reg[31][7]  ( .D(n1546), .CLK(clk), .Q(\regs[31][7] ) );
  DFFX2_LVT \regs_reg[3][12]  ( .D(n2447), .CLK(clk), .Q(\regs[3][12] ) );
  DFFX2_LVT \regs_reg[12][12]  ( .D(n2159), .CLK(clk), .Q(\regs[12][12] ) );
  DFFX2_LVT \regs_reg[14][8]  ( .D(n2091), .CLK(clk), .Q(\regs[14][8] ) );
  DFFX2_LVT \regs_reg[5][2]  ( .D(n2373), .CLK(clk), .Q(\regs[5][2] ) );
  DFFX2_LVT \regs_reg[26][27]  ( .D(n1726), .CLK(clk), .Q(\regs[26][27] ) );
  DFFX2_LVT \regs_reg[31][16]  ( .D(n1555), .CLK(clk), .Q(\regs[31][16] ) );
  DFFX2_LVT \regs_reg[1][2]  ( .D(n2501), .CLK(clk), .Q(\regs[1][2] ) );
  DFFX2_LVT \regs_reg[30][2]  ( .D(n1573), .CLK(clk), .Q(\regs[30][2] ) );
  DFFX2_LVT \regs_reg[25][11]  ( .D(n1742), .CLK(clk), .Q(\regs[25][11] ) );
  DFFX2_LVT \regs_reg[14][21]  ( .D(n2104), .CLK(clk), .Q(\regs[14][21] ) );
  DFFX2_LVT \regs_reg[23][25]  ( .D(n1820), .CLK(clk), .Q(\regs[23][25] ) );
  DFFX2_LVT \regs_reg[9][12]  ( .D(n2255), .CLK(clk), .Q(\regs[9][12] ) );
  DFFX2_LVT \regs_reg[6][11]  ( .D(n2350), .CLK(clk), .Q(\regs[6][11] ) );
  DFFX2_LVT \regs_reg[10][27]  ( .D(n2238), .CLK(clk), .Q(\regs[10][27] ) );
  DFFX2_LVT \regs_reg[19][16]  ( .D(n1939), .CLK(clk), .Q(\regs[19][16] ) );
  DFFX2_LVT \regs_reg[7][16]  ( .D(n2323), .CLK(clk), .Q(\regs[7][16] ) );
  DFFX2_LVT \regs_reg[6][9]  ( .D(n2348), .CLK(clk), .Q(\regs[6][9] ) );
  DFFX2_LVT \regs_reg[9][4]  ( .D(n2247), .CLK(clk), .Q(\regs[9][4] ) );
  DFFX2_LVT \regs_reg[28][16]  ( .D(n1651), .CLK(clk), .Q(\regs[28][16] ) );
  DFFX2_LVT \regs_reg[30][6]  ( .D(n1577), .CLK(clk), .Q(\regs[30][6] ) );
  DFFX2_LVT \regs_reg[1][12]  ( .D(n2511), .CLK(clk), .Q(\regs[1][12] ) );
  DFFX2_LVT \regs_reg[9][30]  ( .D(n2273), .CLK(clk), .Q(\regs[9][30] ) );
  DFFX2_LVT \regs_reg[29][11]  ( .D(n1614), .CLK(clk), .Q(\regs[29][11] ) );
  DFFX2_LVT \regs_reg[4][9]  ( .D(n2412), .CLK(clk), .Q(\regs[4][9] ) );
  DFFX2_LVT \regs_reg[1][30]  ( .D(n2529), .CLK(clk), .Q(\regs[1][30] ) );
  DFFX2_LVT \regs_reg[8][6]  ( .D(n2281), .CLK(clk), .Q(\regs[8][6] ) );
  NBUFFX8_LVT U48 ( .A(n3115), .Y(n3309) );
  NBUFFX8_LVT U303 ( .A(n3096), .Y(n3409) );
  DFFX2_LVT \regs_reg[26][14]  ( .D(n1713), .CLK(clk), .Q(\regs[26][14] ) );
  DFFX2_LVT \regs_reg[29][14]  ( .D(n1617), .CLK(clk), .Q(\regs[29][14] ) );
  DFFX2_LVT \regs_reg[6][29]  ( .D(n2368), .CLK(clk), .Q(\regs[6][29] ) );
  DFFX2_LVT \regs_reg[1][22]  ( .D(n2521), .CLK(clk), .Q(\regs[1][22] ) );
  INVX4_LVT U128 ( .A(n3348), .Y(n3349) );
  DFFX2_LVT \regs_reg[3][29]  ( .D(n2464), .CLK(clk), .Q(\regs[3][29] ) );
  DFFX2_LVT \regs_reg[22][7]  ( .D(n1834), .CLK(clk), .Q(\regs[22][7] ) );
  DFFX2_LVT \regs_reg[23][28]  ( .D(n1823), .CLK(clk), .Q(\regs[23][28] ) );
  DFFX2_LVT \regs_reg[25][10]  ( .D(n1741), .CLK(clk), .Q(\regs[25][10] ) );
  DFFX2_LVT \regs_reg[5][13]  ( .D(n2384), .CLK(clk), .Q(\regs[5][13] ) );
  DFFX2_LVT \regs_reg[3][28]  ( .D(n2463), .CLK(clk), .Q(\regs[3][28] ) );
  DFFX2_LVT \regs_reg[9][29]  ( .D(n2272), .CLK(clk), .Q(\regs[9][29] ) );
  DFFX2_LVT \regs_reg[10][13]  ( .D(n2224), .CLK(clk), .Q(\regs[10][13] ) );
  DFFX2_LVT \regs_reg[5][23]  ( .D(n2394), .CLK(clk), .Q(\regs[5][23] ) );
  DFFX2_LVT \regs_reg[28][29]  ( .D(n1664), .CLK(clk), .Q(\regs[28][29] ) );
  DFFX2_LVT \regs_reg[12][19]  ( .D(n2166), .CLK(clk), .Q(\regs[12][19] ) );
  DFFX2_LVT \regs_reg[19][23]  ( .D(n1946), .CLK(clk), .Q(\regs[19][23] ) );
  DFFX2_LVT \regs_reg[19][9]  ( .D(n1932), .CLK(clk), .Q(\regs[19][9] ) );
  INVX2_LVT U489 ( .A(n3421), .Y(n3422) );
  DFFX2_LVT \regs_reg[27][14]  ( .D(n1681), .CLK(clk), .Q(\regs[27][14] ) );
  DFFX2_LVT \regs_reg[26][18]  ( .D(n1717), .CLK(clk), .Q(\regs[26][18] ) );
  DFFX2_LVT \regs_reg[5][29]  ( .D(n2400), .CLK(clk), .Q(\regs[5][29] ) );
  DFFX2_LVT \regs_reg[22][18]  ( .D(n1845), .CLK(clk), .Q(\regs[22][18] ) );
  DFFX2_LVT \regs_reg[1][28]  ( .D(n2527), .CLK(clk), .Q(\regs[1][28] ) );
  DFFX2_LVT \regs_reg[5][26]  ( .D(n2397), .CLK(clk), .Q(\regs[5][26] ) );
  DFFX2_LVT \regs_reg[23][9]  ( .D(n1804), .CLK(clk), .Q(\regs[23][9] ) );
  DFFX2_LVT \regs_reg[19][10]  ( .D(n1933), .CLK(clk), .Q(\regs[19][10] ) );
  DFFX2_LVT \regs_reg[12][28]  ( .D(n2175), .CLK(clk), .Q(\regs[12][28] ) );
  DFFX2_LVT \regs_reg[8][10]  ( .D(n2285), .CLK(clk), .Q(\regs[8][10] ) );
  DFFX2_LVT \regs_reg[20][13]  ( .D(n1904), .CLK(clk), .Q(\regs[20][13] ) );
  DFFX2_LVT \regs_reg[26][19]  ( .D(n1718), .CLK(clk), .Q(\regs[26][19] ) );
  DFFX2_LVT \regs_reg[23][4]  ( .D(n1799), .CLK(clk), .Q(\regs[23][4] ) );
  DFFX2_LVT \regs_reg[17][28]  ( .D(n2015), .CLK(clk), .Q(\regs[17][28] ) );
  DFFX2_LVT \regs_reg[17][23]  ( .D(n2010), .CLK(clk), .Q(\regs[17][23] ) );
  DFFX2_LVT \regs_reg[1][10]  ( .D(n2509), .CLK(clk), .Q(\regs[1][10] ) );
  DFFX2_LVT \regs_reg[11][7]  ( .D(n2186), .CLK(clk), .Q(\regs[11][7] ) );
  DFFX2_LVT \regs_reg[14][5]  ( .D(n2088), .CLK(clk), .Q(\regs[14][5] ) );
  DFFX2_LVT \regs_reg[3][10]  ( .D(n2445), .CLK(clk), .Q(\regs[3][10] ) );
  DFFX2_LVT \regs_reg[29][29]  ( .D(n1632), .CLK(clk), .Q(\regs[29][29] ) );
  DFFX2_LVT \regs_reg[7][10]  ( .D(n2317), .CLK(clk), .Q(\regs[7][10] ) );
  DFFX2_LVT \regs_reg[25][14]  ( .D(n1745), .CLK(clk), .Q(\regs[25][14] ) );
  DFFX2_LVT \regs_reg[18][19]  ( .D(n1974), .CLK(clk), .Q(\regs[18][19] ) );
  DFFX2_LVT \regs_reg[1][19]  ( .D(n2518), .CLK(clk), .Q(\regs[1][19] ) );
  DFFX2_LVT \regs_reg[15][10]  ( .D(n2061), .CLK(clk), .Q(\regs[15][10] ) );
  DFFX2_LVT \regs_reg[22][22]  ( .D(n1849), .CLK(clk), .Q(\regs[22][22] ) );
  DFFX2_LVT \regs_reg[4][29]  ( .D(n2432), .CLK(clk), .Q(\regs[4][29] ) );
  DFFX2_LVT \regs_reg[21][23]  ( .D(n1882), .CLK(clk), .Q(\regs[21][23] ) );
  DFFX2_LVT \regs_reg[31][4]  ( .D(n1543), .CLK(clk), .Q(\regs[31][4] ) );
  DFFX2_LVT \regs_reg[21][22]  ( .D(n1881), .CLK(clk), .Q(\regs[21][22] ) );
  DFFX2_LVT \regs_reg[2][22]  ( .D(n2489), .CLK(clk), .Q(\regs[2][22] ) );
  DFFX2_LVT \regs_reg[24][17]  ( .D(n1780), .CLK(clk), .Q(\regs[24][17] ) );
  DFFX2_LVT \regs_reg[24][18]  ( .D(n1781), .CLK(clk), .Q(\regs[24][18] ) );
  DFFX2_LVT \regs_reg[20][10]  ( .D(n1901), .CLK(clk), .Q(\regs[20][10] ) );
  DFFX2_LVT \regs_reg[2][13]  ( .D(n2480), .CLK(clk), .Q(\regs[2][13] ) );
  DFFX2_LVT \regs_reg[25][29]  ( .D(n1760), .CLK(clk), .Q(\regs[25][29] ) );
  DFFX2_LVT \regs_reg[30][18]  ( .D(n1589), .CLK(clk), .Q(\regs[30][18] ) );
  DFFX2_LVT \regs_reg[25][8]  ( .D(n1739), .CLK(clk), .Q(\regs[25][8] ) );
  DFFX2_LVT \regs_reg[18][14]  ( .D(n1969), .CLK(clk), .Q(\regs[18][14] ) );
  DFFX2_LVT \regs_reg[25][22]  ( .D(n1753), .CLK(clk), .Q(\regs[25][22] ) );
  DFFX2_LVT \regs_reg[11][6]  ( .D(n2185), .CLK(clk), .Q(\regs[11][6] ) );
  DFFX2_LVT \regs_reg[20][27]  ( .D(n1918), .CLK(clk), .Q(\regs[20][27] ) );
  DFFX2_LVT \regs_reg[18][9]  ( .D(n1964), .CLK(clk), .Q(\regs[18][9] ) );
  DFFX2_LVT \regs_reg[25][16]  ( .D(n1747), .CLK(clk), .Q(\regs[25][16] ) );
  DFFX2_LVT \regs_reg[2][2]  ( .D(n2469), .CLK(clk), .Q(\regs[2][2] ) );
  DFFX2_LVT \regs_reg[22][9]  ( .D(n1836), .CLK(clk), .Q(\regs[22][9] ) );
  DFFX2_LVT \regs_reg[30][23]  ( .D(n1594), .CLK(clk), .Q(\regs[30][23] ) );
  DFFX2_LVT \regs_reg[3][6]  ( .D(n2441), .CLK(clk), .Q(\regs[3][6] ) );
  DFFX2_LVT \regs_reg[13][21]  ( .D(n2136), .CLK(clk), .Q(\regs[13][21] ) );
  DFFX2_LVT \regs_reg[2][12]  ( .D(n2479), .CLK(clk), .Q(\regs[2][12] ) );
  DFFX2_LVT \regs_reg[26][24]  ( .D(n1723), .CLK(clk), .Q(\regs[26][24] ) );
  DFFX2_LVT \regs_reg[14][17]  ( .D(n2100), .CLK(clk), .Q(\regs[14][17] ) );
  DFFX2_LVT \regs_reg[23][10]  ( .D(n1805), .CLK(clk), .Q(\regs[23][10] ) );
  DFFX2_LVT \regs_reg[25][24]  ( .D(n1755), .CLK(clk), .Q(\regs[25][24] ) );
  DFFX2_LVT \regs_reg[26][20]  ( .D(n1719), .CLK(clk), .Q(\regs[26][20] ) );
  DFFX2_LVT \regs_reg[16][4]  ( .D(n2023), .CLK(clk), .Q(\regs[16][4] ) );
  DFFX2_LVT \regs_reg[21][17]  ( .D(n1876), .CLK(clk), .Q(\regs[21][17] ) );
  DFFX2_LVT \regs_reg[8][26]  ( .D(n2301), .CLK(clk), .Q(\regs[8][26] ) );
  DFFX2_LVT \regs_reg[8][14]  ( .D(n2289), .CLK(clk), .Q(\regs[8][14] ) );
  DFFX2_LVT \regs_reg[8][11]  ( .D(n2286), .CLK(clk), .Q(\regs[8][11] ) );
  DFFX2_LVT \regs_reg[4][19]  ( .D(n2422), .CLK(clk), .Q(\regs[4][19] ) );
  DFFX2_LVT \regs_reg[28][19]  ( .D(n1654), .CLK(clk), .Q(\regs[28][19] ) );
  INVX4_LVT U98 ( .A(n3331), .Y(n3332) );
  DFFX2_LVT \regs_reg[10][18]  ( .D(n2229), .CLK(clk), .Q(\regs[10][18] ) );
  DFFX2_LVT \regs_reg[23][18]  ( .D(n1813), .CLK(clk), .Q(\regs[23][18] ) );
  INVX4_LVT U435 ( .A(n3417), .Y(n3418) );
  DFFX2_LVT \regs_reg[29][31]  ( .D(n1634), .CLK(clk), .Q(\regs[29][31] ) );
  DFFX2_LVT \regs_reg[25][23]  ( .D(n1754), .CLK(clk), .Q(\regs[25][23] ) );
  INVX4_LVT U523 ( .A(n3424), .Y(n3425) );
  DFFX2_LVT \regs_reg[28][23]  ( .D(n1658), .CLK(clk), .Q(\regs[28][23] ) );
  DFFX2_LVT \regs_reg[17][20]  ( .D(n2007), .CLK(clk), .Q(\regs[17][20] ) );
  DFFX2_LVT \regs_reg[3][31]  ( .D(n2466), .CLK(clk), .Q(\regs[3][31] ) );
  DFFX2_LVT \regs_reg[23][20]  ( .D(n1815), .CLK(clk), .Q(\regs[23][20] ) );
  DFFX2_LVT \regs_reg[22][20]  ( .D(n1847), .CLK(clk), .Q(\regs[22][20] ) );
  DFFX2_LVT \regs_reg[8][17]  ( .D(n2292), .CLK(clk), .Q(\regs[8][17] ) );
  DFFX2_LVT \regs_reg[8][8]  ( .D(n2283), .CLK(clk), .Q(\regs[8][8] ) );
  DFFX2_LVT \regs_reg[13][6]  ( .D(n2121), .CLK(clk), .Q(\regs[13][6] ) );
  DFFX2_LVT \regs_reg[15][28]  ( .D(n2079), .CLK(clk), .Q(\regs[15][28] ) );
  DFFX2_LVT \regs_reg[5][16]  ( .D(n2387), .CLK(clk), .Q(\regs[5][16] ) );
  DFFX2_LVT \regs_reg[27][27]  ( .D(n1694), .CLK(clk), .Q(\regs[27][27] ) );
  DFFX2_LVT \regs_reg[29][23]  ( .D(n1626), .CLK(clk), .Q(\regs[29][23] ) );
  DFFX2_LVT \regs_reg[22][25]  ( .D(n1852), .CLK(clk), .Q(\regs[22][25] ) );
  DFFX2_LVT \regs_reg[26][22]  ( .D(n1721), .CLK(clk), .Q(\regs[26][22] ) );
  DFFX2_LVT \regs_reg[30][24]  ( .D(n1595), .CLK(clk), .Q(\regs[30][24] ) );
  DFFX2_LVT \regs_reg[30][25]  ( .D(n1596), .CLK(clk), .Q(\regs[30][25] ) );
  DFFX2_LVT \regs_reg[1][3]  ( .D(n2502), .CLK(clk), .Q(\regs[1][3] ) );
  DFFX2_LVT \regs_reg[15][5]  ( .D(n2056), .CLK(clk), .Q(\regs[15][5] ) );
  DFFX2_LVT \regs_reg[8][7]  ( .D(n2282), .CLK(clk), .Q(\regs[8][7] ) );
  DFFX2_LVT \regs_reg[25][5]  ( .D(n1736), .CLK(clk), .Q(\regs[25][5] ) );
  DFFX2_LVT \regs_reg[25][7]  ( .D(n1738), .CLK(clk), .Q(\regs[25][7] ) );
  DFFX2_LVT \regs_reg[23][8]  ( .D(n1803), .CLK(clk), .Q(\regs[23][8] ) );
  DFFX2_LVT \regs_reg[3][14]  ( .D(n2449), .CLK(clk), .Q(\regs[3][14] ) );
  DFFX2_LVT \regs_reg[5][6]  ( .D(n2377), .CLK(clk), .Q(\regs[5][6] ) );
  DFFX2_LVT \regs_reg[11][9]  ( .D(n2188), .CLK(clk), .Q(\regs[11][9] ) );
  DFFX2_LVT \regs_reg[28][10]  ( .D(n1645), .CLK(clk), .Q(\regs[28][10] ) );
  DFFX2_LVT \regs_reg[25][6]  ( .D(n1737), .CLK(clk), .Q(\regs[25][6] ) );
  DFFX2_LVT \regs_reg[4][4]  ( .D(n2407), .CLK(clk), .Q(\regs[4][4] ) );
  DFFX2_LVT \regs_reg[29][18]  ( .D(n1621), .CLK(clk), .Q(\regs[29][18] ) );
  DFFX2_LVT \regs_reg[22][19]  ( .D(n1846), .CLK(clk), .Q(\regs[22][19] ) );
  DFFX2_LVT \regs_reg[18][30]  ( .D(n1985), .CLK(clk), .Q(\regs[18][30] ) );
  DFFX2_LVT \regs_reg[28][12]  ( .D(n1647), .CLK(clk), .Q(\regs[28][12] ) );
  DFFX2_LVT \regs_reg[29][19]  ( .D(n1622), .CLK(clk), .Q(\regs[29][19] ) );
  INVX4_LVT U166 ( .A(n3363), .Y(n3366) );
  DFFX2_LVT \regs_reg[27][22]  ( .D(n1689), .CLK(clk), .Q(\regs[27][22] ) );
  DFFX2_LVT \regs_reg[21][20]  ( .D(n1879), .CLK(clk), .Q(\regs[21][20] ) );
  DFFX2_LVT \regs_reg[21][24]  ( .D(n1883), .CLK(clk), .Q(\regs[21][24] ) );
  DFFX2_LVT \regs_reg[8][5]  ( .D(n2280), .CLK(clk), .Q(\regs[8][5] ) );
  DFFX2_LVT \regs_reg[20][19]  ( .D(n1910), .CLK(clk), .Q(\regs[20][19] ) );
  DFFX2_LVT \regs_reg[29][20]  ( .D(n1623), .CLK(clk), .Q(\regs[29][20] ) );
  DFFX2_LVT \regs_reg[25][18]  ( .D(n1749), .CLK(clk), .Q(\regs[25][18] ) );
  DFFX2_LVT \regs_reg[26][3]  ( .D(n1702), .CLK(clk), .Q(\regs[26][3] ) );
  DFFX2_LVT \regs_reg[19][15]  ( .D(n1938), .CLK(clk), .Q(\regs[19][15] ) );
  DFFX2_LVT \regs_reg[18][5]  ( .D(n1960), .CLK(clk), .Q(\regs[18][5] ) );
  DFFX2_LVT \regs_reg[6][14]  ( .D(n2353), .CLK(clk), .Q(\regs[6][14] ) );
  NBUFFX8_LVT U127 ( .A(n3068), .Y(n3348) );
  NAND3X2_LVT U2249 ( .A1(n3470), .A2(n3202), .A3(n2992), .Y(n2974) );
  DFFX2_LVT \regs_reg[7][3]  ( .D(n2310), .CLK(clk), .Q(\regs[7][3] ) );
  DFFX2_LVT \regs_reg[5][5]  ( .D(n2376), .CLK(clk), .Q(\regs[5][5] ) );
  DFFX2_LVT \regs_reg[28][13]  ( .D(n1648), .CLK(clk), .Q(\regs[28][13] ) );
  DFFX2_LVT \regs_reg[12][26]  ( .D(n2173), .CLK(clk), .Q(\regs[12][26] ) );
  DFFX2_LVT \regs_reg[28][24]  ( .D(n1659), .CLK(clk), .Q(\regs[28][24] ) );
  DFFX2_LVT \regs_reg[30][26]  ( .D(n1597), .CLK(clk), .Q(\regs[30][26] ) );
  DFFX2_LVT \regs_reg[31][24]  ( .D(n1563), .CLK(clk), .Q(\regs[31][24] ) );
  NAND3X2_LVT U2661 ( .A1(n3470), .A2(n3255), .A3(n3067), .Y(n3068) );
  DFFX2_LVT \regs_reg[24][4]  ( .D(n1767), .CLK(clk), .Q(\regs[24][4] ) );
  NBUFFX8_LVT U156 ( .A(n2993), .Y(n3363) );
  NAND3X2_LVT U2331 ( .A1(n3470), .A2(n2992), .A3(n3255), .Y(n2993) );
  NBUFFX4_LVT U130 ( .A(n1027), .Y(n3481) );
  NBUFFX4_LVT U161 ( .A(n969), .Y(n3475) );
  NBUFFX4_LVT U193 ( .A(waddr[2]), .Y(n3470) );
  NBUFFX4_LVT U995 ( .A(wdata[20]), .Y(n3469) );
  NBUFFX4_LVT U1021 ( .A(wdata[29]), .Y(n3453) );
  NBUFFX4_LVT U1023 ( .A(n148), .Y(n3454) );
  NBUFFX4_LVT U1024 ( .A(n135), .Y(n3455) );
  NBUFFX4_LVT U1025 ( .A(n26), .Y(n3456) );
  NBUFFX4_LVT U1032 ( .A(n56), .Y(n3457) );
  NBUFFX4_LVT U1042 ( .A(n52), .Y(n3458) );
  NBUFFX4_LVT U1043 ( .A(n30), .Y(n3459) );
  NBUFFX4_LVT U1045 ( .A(n120), .Y(n3460) );
  NBUFFX4_LVT U1046 ( .A(n37), .Y(n3461) );
  NBUFFX4_LVT U1050 ( .A(n110), .Y(n3462) );
  NBUFFX4_LVT U1051 ( .A(n40), .Y(n3463) );
  NBUFFX4_LVT U1055 ( .A(n24), .Y(n3464) );
  NBUFFX4_LVT U1056 ( .A(n122), .Y(n3465) );
  NBUFFX4_LVT U1060 ( .A(n11), .Y(n3466) );
  NBUFFX4_LVT U1061 ( .A(n63), .Y(n3467) );
  NBUFFX4_LVT U1063 ( .A(n50), .Y(n3468) );
  NBUFFX4_LVT U1064 ( .A(n9), .Y(n3471) );
  NBUFFX4_LVT U1069 ( .A(n38), .Y(n3472) );
  NBUFFX4_LVT U1070 ( .A(n21), .Y(n3473) );
  NBUFFX4_LVT U1072 ( .A(n58), .Y(n3474) );
  NBUFFX4_LVT U1073 ( .A(n25), .Y(n3476) );
  NBUFFX4_LVT U1077 ( .A(n54), .Y(n3477) );
  NBUFFX4_LVT U1078 ( .A(n61), .Y(n3478) );
  NBUFFX4_LVT U1083 ( .A(n28), .Y(n3479) );
  NBUFFX4_LVT U1084 ( .A(n42), .Y(n3480) );
  NBUFFX4_LVT U1087 ( .A(n29), .Y(n3482) );
  NBUFFX8_LVT U1088 ( .A(n3492), .Y(n3483) );
  NBUFFX4_LVT U1091 ( .A(n23), .Y(n3484) );
  NBUFFX4_LVT U1092 ( .A(n43), .Y(n3485) );
  NBUFFX8_LVT U1095 ( .A(wdata[31]), .Y(n3486) );
  NBUFFX4_LVT U1096 ( .A(n65), .Y(n3487) );
  NBUFFX8_LVT U1100 ( .A(wdata[22]), .Y(n3494) );
  NBUFFX8_LVT U1101 ( .A(wdata[23]), .Y(n3497) );
  NBUFFX8_LVT U1103 ( .A(wdata[24]), .Y(n3493) );
  NBUFFX8_LVT U1104 ( .A(wdata[19]), .Y(n3496) );
  NBUFFX8_LVT U1107 ( .A(wdata[18]), .Y(n3491) );
  NBUFFX8_LVT U1108 ( .A(n3453), .Y(n3501) );
  NBUFFX8_LVT U1111 ( .A(wdata[13]), .Y(n3502) );
  NBUFFX8_LVT U1112 ( .A(wdata[14]), .Y(n3498) );
  NBUFFX8_LVT U1116 ( .A(wdata[15]), .Y(n3495) );
  NBUFFX8_LVT U1117 ( .A(wdata[10]), .Y(n3499) );
  NBUFFX8_LVT U1119 ( .A(wdata[28]), .Y(n3500) );
  NBUFFX8_LVT U1120 ( .A(wdata[26]), .Y(n3503) );
  NBUFFX4_LVT U1123 ( .A(n39), .Y(n3488) );
  NBUFFX4_LVT U1124 ( .A(n36), .Y(n3489) );
  NBUFFX4_LVT U1126 ( .A(n44), .Y(n3490) );
  NBUFFX4_LVT U1127 ( .A(n3469), .Y(n3492) );
endmodule


module pipe_id_ex ( clk, rst, id_aluop, id_alusel, id_opv1, id_opv2, 
        id_reg_waddr, id_we, stall, id_link_addr, id_mem_offset, ex_aluop, 
        ex_alusel, ex_opv1, ex_opv2, ex_reg_waddr, ex_we, ex_link_addr, 
        ex_mem_offset );
  input [7:0] id_aluop;
  input [2:0] id_alusel;
  input [31:0] id_opv1;
  input [31:0] id_opv2;
  input [4:0] id_reg_waddr;
  input [5:0] stall;
  input [31:0] id_link_addr;
  input [31:0] id_mem_offset;
  output [7:0] ex_aluop;
  output [2:0] ex_alusel;
  output [31:0] ex_opv1;
  output [31:0] ex_opv2;
  output [4:0] ex_reg_waddr;
  output [31:0] ex_link_addr;
  output [31:0] ex_mem_offset;
  input clk, rst, id_we;
  output ex_we;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n173, n175, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195;

  DFFX1_LVT \ex_link_addr_reg[30]  ( .D(n144), .CLK(clk), .Q(ex_link_addr[30])
         );
  DFFX1_LVT \ex_link_addr_reg[31]  ( .D(n145), .CLK(clk), .Q(ex_link_addr[31])
         );
  DFFX1_LVT \ex_link_addr_reg[17]  ( .D(n131), .CLK(clk), .Q(ex_link_addr[17])
         );
  DFFX1_LVT \ex_link_addr_reg[22]  ( .D(n136), .CLK(clk), .Q(ex_link_addr[22])
         );
  DFFX1_LVT \ex_link_addr_reg[9]  ( .D(n123), .CLK(clk), .Q(ex_link_addr[9])
         );
  DFFX1_LVT \ex_link_addr_reg[0]  ( .D(n114), .CLK(clk), .Q(ex_link_addr[0])
         );
  DFFX1_LVT \ex_link_addr_reg[6]  ( .D(n120), .CLK(clk), .Q(ex_link_addr[6])
         );
  DFFX1_LVT \ex_link_addr_reg[14]  ( .D(n128), .CLK(clk), .Q(ex_link_addr[14])
         );
  DFFX1_LVT \ex_link_addr_reg[28]  ( .D(n142), .CLK(clk), .Q(ex_link_addr[28])
         );
  DFFX1_LVT \ex_link_addr_reg[15]  ( .D(n129), .CLK(clk), .Q(ex_link_addr[15])
         );
  DFFX1_LVT \ex_link_addr_reg[16]  ( .D(n130), .CLK(clk), .Q(ex_link_addr[16])
         );
  DFFX1_LVT \ex_link_addr_reg[4]  ( .D(n118), .CLK(clk), .Q(ex_link_addr[4])
         );
  DFFX1_LVT \ex_link_addr_reg[27]  ( .D(n141), .CLK(clk), .Q(ex_link_addr[27])
         );
  DFFX1_LVT \ex_link_addr_reg[26]  ( .D(n140), .CLK(clk), .Q(ex_link_addr[26])
         );
  DFFX1_LVT \ex_mem_offset_reg[30]  ( .D(n112), .CLK(clk), .Q(
        ex_mem_offset[30]) );
  DFFX1_LVT \ex_link_addr_reg[8]  ( .D(n122), .CLK(clk), .Q(ex_link_addr[8])
         );
  DFFX1_LVT \ex_link_addr_reg[7]  ( .D(n121), .CLK(clk), .Q(ex_link_addr[7])
         );
  DFFX1_LVT \ex_link_addr_reg[5]  ( .D(n119), .CLK(clk), .Q(ex_link_addr[5])
         );
  DFFX1_LVT \ex_link_addr_reg[24]  ( .D(n138), .CLK(clk), .Q(ex_link_addr[24])
         );
  DFFX1_LVT \ex_link_addr_reg[19]  ( .D(n133), .CLK(clk), .Q(ex_link_addr[19])
         );
  DFFX1_LVT \ex_link_addr_reg[23]  ( .D(n137), .CLK(clk), .Q(ex_link_addr[23])
         );
  DFFX1_LVT \ex_link_addr_reg[11]  ( .D(n125), .CLK(clk), .Q(ex_link_addr[11])
         );
  DFFX1_LVT \ex_link_addr_reg[3]  ( .D(n117), .CLK(clk), .Q(ex_link_addr[3])
         );
  DFFX1_LVT \ex_link_addr_reg[20]  ( .D(n134), .CLK(clk), .Q(ex_link_addr[20])
         );
  DFFX1_LVT \ex_mem_offset_reg[31]  ( .D(n113), .CLK(clk), .Q(
        ex_mem_offset[31]) );
  DFFX1_LVT \ex_link_addr_reg[18]  ( .D(n132), .CLK(clk), .Q(ex_link_addr[18])
         );
  DFFX1_LVT \ex_link_addr_reg[29]  ( .D(n143), .CLK(clk), .Q(ex_link_addr[29])
         );
  DFFX1_LVT \ex_link_addr_reg[1]  ( .D(n115), .CLK(clk), .Q(ex_link_addr[1])
         );
  DFFX1_LVT \ex_link_addr_reg[2]  ( .D(n116), .CLK(clk), .Q(ex_link_addr[2])
         );
  DFFX1_LVT \ex_link_addr_reg[13]  ( .D(n127), .CLK(clk), .Q(ex_link_addr[13])
         );
  DFFX1_LVT \ex_link_addr_reg[12]  ( .D(n126), .CLK(clk), .Q(ex_link_addr[12])
         );
  DFFX1_LVT \ex_link_addr_reg[21]  ( .D(n135), .CLK(clk), .Q(ex_link_addr[21])
         );
  DFFX1_LVT \ex_link_addr_reg[25]  ( .D(n139), .CLK(clk), .Q(ex_link_addr[25])
         );
  DFFX1_LVT \ex_link_addr_reg[10]  ( .D(n124), .CLK(clk), .Q(ex_link_addr[10])
         );
  DFFX1_LVT \ex_mem_offset_reg[29]  ( .D(n111), .CLK(clk), .Q(
        ex_mem_offset[29]) );
  DFFX1_LVT \ex_mem_offset_reg[28]  ( .D(n110), .CLK(clk), .Q(
        ex_mem_offset[28]) );
  DFFX1_LVT \ex_opv2_reg[31]  ( .D(n41), .CLK(clk), .Q(ex_opv2[31]) );
  DFFX1_LVT \ex_mem_offset_reg[27]  ( .D(n109), .CLK(clk), .Q(
        ex_mem_offset[27]) );
  DFFX1_LVT \ex_opv2_reg[30]  ( .D(n40), .CLK(clk), .Q(ex_opv2[30]) );
  DFFX1_LVT \ex_mem_offset_reg[26]  ( .D(n108), .CLK(clk), .Q(
        ex_mem_offset[26]) );
  DFFX1_LVT \ex_opv2_reg[29]  ( .D(n39), .CLK(clk), .Q(ex_opv2[29]) );
  DFFX1_LVT \ex_opv2_reg[28]  ( .D(n38), .CLK(clk), .Q(ex_opv2[28]) );
  DFFX1_LVT \ex_mem_offset_reg[25]  ( .D(n107), .CLK(clk), .Q(
        ex_mem_offset[25]) );
  DFFX1_LVT \ex_mem_offset_reg[24]  ( .D(n106), .CLK(clk), .Q(
        ex_mem_offset[24]) );
  DFFX1_LVT \ex_mem_offset_reg[23]  ( .D(n105), .CLK(clk), .Q(
        ex_mem_offset[23]) );
  DFFX1_LVT \ex_opv2_reg[26]  ( .D(n36), .CLK(clk), .Q(ex_opv2[26]) );
  DFFX1_LVT \ex_opv2_reg[25]  ( .D(n35), .CLK(clk), .Q(ex_opv2[25]) );
  DFFX1_LVT \ex_opv2_reg[27]  ( .D(n37), .CLK(clk), .Q(ex_opv2[27]) );
  DFFX1_LVT \ex_mem_offset_reg[22]  ( .D(n104), .CLK(clk), .Q(
        ex_mem_offset[22]) );
  DFFX1_LVT \ex_opv2_reg[24]  ( .D(n34), .CLK(clk), .Q(ex_opv2[24]) );
  DFFX1_LVT \ex_mem_offset_reg[21]  ( .D(n103), .CLK(clk), .Q(
        ex_mem_offset[21]) );
  DFFX1_LVT \ex_alusel_reg[1]  ( .D(n75), .CLK(clk), .Q(ex_alusel[1]) );
  DFFX1_LVT \ex_alusel_reg[0]  ( .D(n74), .CLK(clk), .Q(ex_alusel[0]) );
  DFFX1_LVT \ex_opv2_reg[23]  ( .D(n33), .CLK(clk), .Q(ex_opv2[23]) );
  DFFX1_LVT \ex_alusel_reg[2]  ( .D(n76), .CLK(clk), .Q(ex_alusel[2]) );
  DFFX1_LVT \ex_mem_offset_reg[20]  ( .D(n102), .CLK(clk), .Q(
        ex_mem_offset[20]) );
  DFFX1_LVT \ex_opv2_reg[22]  ( .D(n32), .CLK(clk), .Q(ex_opv2[22]) );
  DFFX1_LVT \ex_mem_offset_reg[19]  ( .D(n101), .CLK(clk), .Q(
        ex_mem_offset[19]) );
  DFFX1_LVT \ex_opv2_reg[21]  ( .D(n31), .CLK(clk), .Q(ex_opv2[21]) );
  DFFX1_LVT \ex_mem_offset_reg[18]  ( .D(n100), .CLK(clk), .Q(
        ex_mem_offset[18]) );
  DFFX1_LVT \ex_aluop_reg[3]  ( .D(n80), .CLK(clk), .Q(ex_aluop[3]) );
  DFFX1_LVT \ex_opv2_reg[20]  ( .D(n30), .CLK(clk), .Q(ex_opv2[20]) );
  DFFX1_LVT \ex_reg_waddr_reg[0]  ( .D(n5), .CLK(clk), .Q(ex_reg_waddr[0]) );
  DFFX1_LVT \ex_reg_waddr_reg[1]  ( .D(n6), .CLK(clk), .Q(ex_reg_waddr[1]) );
  DFFX1_LVT \ex_reg_waddr_reg[2]  ( .D(n7), .CLK(clk), .Q(ex_reg_waddr[2]) );
  DFFX1_LVT \ex_reg_waddr_reg[4]  ( .D(n9), .CLK(clk), .Q(ex_reg_waddr[4]) );
  DFFX1_LVT \ex_reg_waddr_reg[3]  ( .D(n8), .CLK(clk), .Q(ex_reg_waddr[3]) );
  DFFX1_LVT \ex_mem_offset_reg[17]  ( .D(n99), .CLK(clk), .Q(ex_mem_offset[17]) );
  DFFX1_LVT \ex_opv2_reg[19]  ( .D(n29), .CLK(clk), .Q(ex_opv2[19]) );
  DFFX1_LVT \ex_mem_offset_reg[16]  ( .D(n98), .CLK(clk), .Q(ex_mem_offset[16]) );
  DFFX1_LVT \ex_opv2_reg[18]  ( .D(n28), .CLK(clk), .Q(ex_opv2[18]) );
  DFFX1_LVT \ex_mem_offset_reg[15]  ( .D(n97), .CLK(clk), .Q(ex_mem_offset[15]) );
  DFFX1_LVT \ex_opv2_reg[17]  ( .D(n27), .CLK(clk), .Q(ex_opv2[17]) );
  DFFX1_LVT \ex_mem_offset_reg[14]  ( .D(n96), .CLK(clk), .Q(ex_mem_offset[14]) );
  DFFX1_LVT \ex_opv2_reg[16]  ( .D(n26), .CLK(clk), .Q(ex_opv2[16]) );
  DFFX1_LVT \ex_mem_offset_reg[13]  ( .D(n95), .CLK(clk), .Q(ex_mem_offset[13]) );
  DFFX1_LVT \ex_opv2_reg[15]  ( .D(n25), .CLK(clk), .Q(ex_opv2[15]) );
  DFFX1_LVT \ex_mem_offset_reg[12]  ( .D(n94), .CLK(clk), .Q(ex_mem_offset[12]) );
  DFFX1_LVT \ex_opv2_reg[14]  ( .D(n24), .CLK(clk), .Q(ex_opv2[14]) );
  DFFX1_LVT \ex_mem_offset_reg[11]  ( .D(n93), .CLK(clk), .Q(ex_mem_offset[11]) );
  DFFX1_LVT \ex_opv2_reg[13]  ( .D(n23), .CLK(clk), .Q(ex_opv2[13]) );
  DFFX1_LVT \ex_mem_offset_reg[10]  ( .D(n92), .CLK(clk), .Q(ex_mem_offset[10]) );
  DFFX1_LVT \ex_opv2_reg[12]  ( .D(n22), .CLK(clk), .Q(ex_opv2[12]) );
  DFFX1_LVT \ex_mem_offset_reg[9]  ( .D(n91), .CLK(clk), .Q(ex_mem_offset[9])
         );
  DFFX1_LVT \ex_opv2_reg[11]  ( .D(n21), .CLK(clk), .Q(ex_opv2[11]) );
  DFFX1_LVT \ex_mem_offset_reg[8]  ( .D(n90), .CLK(clk), .Q(ex_mem_offset[8])
         );
  DFFX1_LVT \ex_opv2_reg[10]  ( .D(n20), .CLK(clk), .Q(ex_opv2[10]) );
  DFFX1_LVT \ex_mem_offset_reg[7]  ( .D(n89), .CLK(clk), .Q(ex_mem_offset[7])
         );
  DFFX1_LVT \ex_mem_offset_reg[6]  ( .D(n88), .CLK(clk), .Q(ex_mem_offset[6])
         );
  DFFX1_LVT \ex_opv2_reg[8]  ( .D(n18), .CLK(clk), .Q(ex_opv2[8]) );
  DFFX1_LVT \ex_mem_offset_reg[5]  ( .D(n87), .CLK(clk), .Q(ex_mem_offset[5])
         );
  DFFX1_LVT \ex_opv2_reg[7]  ( .D(n17), .CLK(clk), .Q(ex_opv2[7]) );
  DFFX1_LVT \ex_mem_offset_reg[4]  ( .D(n86), .CLK(clk), .Q(ex_mem_offset[4])
         );
  DFFX1_LVT \ex_opv2_reg[6]  ( .D(n16), .CLK(clk), .Q(ex_opv2[6]) );
  DFFX1_LVT \ex_mem_offset_reg[3]  ( .D(n85), .CLK(clk), .Q(ex_mem_offset[3])
         );
  DFFX1_LVT \ex_opv2_reg[5]  ( .D(n15), .CLK(clk), .Q(ex_opv2[5]) );
  DFFX1_LVT \ex_mem_offset_reg[2]  ( .D(n84), .CLK(clk), .Q(ex_mem_offset[2])
         );
  DFFX1_LVT \ex_opv2_reg[4]  ( .D(n14), .CLK(clk), .Q(ex_opv2[4]) );
  DFFX1_LVT \ex_mem_offset_reg[1]  ( .D(n83), .CLK(clk), .Q(ex_mem_offset[1])
         );
  DFFX1_LVT \ex_opv2_reg[3]  ( .D(n13), .CLK(clk), .Q(ex_opv2[3]) );
  DFFX1_LVT \ex_opv2_reg[2]  ( .D(n12), .CLK(clk), .Q(ex_opv2[2]) );
  DFFX1_LVT \ex_mem_offset_reg[0]  ( .D(n82), .CLK(clk), .Q(ex_mem_offset[0])
         );
  DFFX1_LVT \ex_opv1_reg[0]  ( .D(n42), .CLK(clk), .Q(ex_opv1[0]) );
  DFFX1_LVT \ex_opv2_reg[1]  ( .D(n11), .CLK(clk), .Q(ex_opv2[1]) );
  DFFX1_LVT \ex_opv2_reg[0]  ( .D(n10), .CLK(clk), .Q(ex_opv2[0]) );
  DFFX1_LVT \ex_aluop_reg[0]  ( .D(n77), .CLK(clk), .Q(ex_aluop[0]) );
  AND3X1_LVT U4 ( .A1(stall[2]), .A2(stall[3]), .A3(n185), .Y(n173) );
  NOR2X0_LVT U8 ( .A1(stall[2]), .A2(rst), .Y(n175) );
  AO22X1_LVT U12 ( .A1(n187), .A2(ex_we), .A3(n192), .A4(id_we), .Y(n146) );
  AO22X1_LVT U13 ( .A1(n187), .A2(ex_link_addr[31]), .A3(n192), .A4(
        id_link_addr[31]), .Y(n145) );
  AO22X1_LVT U14 ( .A1(n187), .A2(ex_link_addr[30]), .A3(n192), .A4(
        id_link_addr[30]), .Y(n144) );
  AO22X1_LVT U15 ( .A1(n187), .A2(ex_link_addr[29]), .A3(n192), .A4(
        id_link_addr[29]), .Y(n143) );
  AO22X1_LVT U16 ( .A1(n187), .A2(ex_link_addr[28]), .A3(n192), .A4(
        id_link_addr[28]), .Y(n142) );
  AO22X1_LVT U17 ( .A1(n187), .A2(ex_link_addr[27]), .A3(n192), .A4(
        id_link_addr[27]), .Y(n141) );
  AO22X1_LVT U18 ( .A1(n187), .A2(ex_link_addr[26]), .A3(n192), .A4(
        id_link_addr[26]), .Y(n140) );
  AO22X1_LVT U19 ( .A1(n187), .A2(ex_link_addr[25]), .A3(n192), .A4(
        id_link_addr[25]), .Y(n139) );
  AO22X1_LVT U20 ( .A1(n187), .A2(ex_link_addr[24]), .A3(n192), .A4(
        id_link_addr[24]), .Y(n138) );
  AO22X1_LVT U21 ( .A1(n187), .A2(ex_link_addr[23]), .A3(n192), .A4(
        id_link_addr[23]), .Y(n137) );
  AO22X1_LVT U22 ( .A1(n187), .A2(ex_link_addr[22]), .A3(n192), .A4(
        id_link_addr[22]), .Y(n136) );
  AO22X1_LVT U23 ( .A1(n187), .A2(ex_link_addr[21]), .A3(n192), .A4(
        id_link_addr[21]), .Y(n135) );
  AO22X1_LVT U26 ( .A1(n187), .A2(ex_link_addr[20]), .A3(n192), .A4(
        id_link_addr[20]), .Y(n134) );
  AO22X1_LVT U27 ( .A1(n187), .A2(ex_link_addr[19]), .A3(n192), .A4(
        id_link_addr[19]), .Y(n133) );
  AO22X1_LVT U28 ( .A1(n187), .A2(ex_link_addr[18]), .A3(n192), .A4(
        id_link_addr[18]), .Y(n132) );
  AO22X1_LVT U29 ( .A1(n187), .A2(ex_link_addr[17]), .A3(n192), .A4(
        id_link_addr[17]), .Y(n131) );
  AO22X1_LVT U30 ( .A1(n187), .A2(ex_link_addr[16]), .A3(n192), .A4(
        id_link_addr[16]), .Y(n130) );
  AO22X1_LVT U31 ( .A1(n187), .A2(ex_link_addr[15]), .A3(n192), .A4(
        id_link_addr[15]), .Y(n129) );
  AO22X1_LVT U32 ( .A1(n187), .A2(ex_link_addr[14]), .A3(n192), .A4(
        id_link_addr[14]), .Y(n128) );
  AO22X1_LVT U33 ( .A1(n187), .A2(ex_link_addr[13]), .A3(n192), .A4(
        id_link_addr[13]), .Y(n127) );
  AO22X1_LVT U34 ( .A1(n187), .A2(ex_link_addr[12]), .A3(n192), .A4(
        id_link_addr[12]), .Y(n126) );
  AO22X1_LVT U35 ( .A1(n187), .A2(ex_link_addr[11]), .A3(n192), .A4(
        id_link_addr[11]), .Y(n125) );
  AO22X1_LVT U36 ( .A1(n187), .A2(ex_link_addr[10]), .A3(n192), .A4(
        id_link_addr[10]), .Y(n124) );
  AO22X1_LVT U37 ( .A1(n187), .A2(ex_link_addr[9]), .A3(n192), .A4(
        id_link_addr[9]), .Y(n123) );
  AO22X1_LVT U40 ( .A1(n187), .A2(ex_link_addr[8]), .A3(n192), .A4(
        id_link_addr[8]), .Y(n122) );
  AO22X1_LVT U41 ( .A1(n187), .A2(ex_link_addr[7]), .A3(n192), .A4(
        id_link_addr[7]), .Y(n121) );
  AO22X1_LVT U42 ( .A1(n187), .A2(ex_link_addr[6]), .A3(n192), .A4(
        id_link_addr[6]), .Y(n120) );
  AO22X1_LVT U43 ( .A1(n187), .A2(ex_link_addr[5]), .A3(n192), .A4(
        id_link_addr[5]), .Y(n119) );
  AO22X1_LVT U44 ( .A1(n187), .A2(ex_link_addr[4]), .A3(n192), .A4(
        id_link_addr[4]), .Y(n118) );
  AO22X1_LVT U45 ( .A1(n187), .A2(ex_link_addr[3]), .A3(n192), .A4(
        id_link_addr[3]), .Y(n117) );
  AO22X1_LVT U46 ( .A1(n187), .A2(ex_link_addr[2]), .A3(n192), .A4(
        id_link_addr[2]), .Y(n116) );
  AO22X1_LVT U47 ( .A1(n187), .A2(ex_link_addr[1]), .A3(n192), .A4(
        id_link_addr[1]), .Y(n115) );
  AO22X1_LVT U48 ( .A1(n187), .A2(ex_link_addr[0]), .A3(n192), .A4(
        id_link_addr[0]), .Y(n114) );
  AO22X1_LVT U49 ( .A1(n187), .A2(ex_mem_offset[31]), .A3(n192), .A4(
        id_mem_offset[31]), .Y(n113) );
  AO22X1_LVT U50 ( .A1(n187), .A2(ex_mem_offset[30]), .A3(n192), .A4(
        id_mem_offset[30]), .Y(n112) );
  AO22X1_LVT U51 ( .A1(n187), .A2(ex_mem_offset[29]), .A3(n192), .A4(
        id_mem_offset[29]), .Y(n111) );
  AO22X1_LVT U56 ( .A1(n189), .A2(ex_mem_offset[28]), .A3(n194), .A4(
        id_mem_offset[28]), .Y(n110) );
  AO22X1_LVT U57 ( .A1(n189), .A2(ex_mem_offset[27]), .A3(n194), .A4(
        id_mem_offset[27]), .Y(n109) );
  AO22X1_LVT U58 ( .A1(n189), .A2(ex_mem_offset[26]), .A3(n194), .A4(
        id_mem_offset[26]), .Y(n108) );
  AO22X1_LVT U59 ( .A1(n189), .A2(ex_mem_offset[25]), .A3(n194), .A4(
        id_mem_offset[25]), .Y(n107) );
  AO22X1_LVT U60 ( .A1(n189), .A2(ex_mem_offset[24]), .A3(n194), .A4(
        id_mem_offset[24]), .Y(n106) );
  AO22X1_LVT U61 ( .A1(n189), .A2(ex_mem_offset[23]), .A3(n194), .A4(
        id_mem_offset[23]), .Y(n105) );
  AO22X1_LVT U62 ( .A1(n189), .A2(ex_mem_offset[22]), .A3(n194), .A4(
        id_mem_offset[22]), .Y(n104) );
  AO22X1_LVT U63 ( .A1(n189), .A2(ex_mem_offset[21]), .A3(n194), .A4(
        id_mem_offset[21]), .Y(n103) );
  AO22X1_LVT U64 ( .A1(n189), .A2(ex_mem_offset[20]), .A3(n194), .A4(
        id_mem_offset[20]), .Y(n102) );
  AO22X1_LVT U65 ( .A1(n189), .A2(ex_mem_offset[19]), .A3(n194), .A4(
        id_mem_offset[19]), .Y(n101) );
  AO22X1_LVT U66 ( .A1(n189), .A2(ex_mem_offset[18]), .A3(n194), .A4(
        id_mem_offset[18]), .Y(n100) );
  AO22X1_LVT U67 ( .A1(n189), .A2(ex_mem_offset[17]), .A3(n194), .A4(
        id_mem_offset[17]), .Y(n99) );
  AO22X1_LVT U70 ( .A1(n189), .A2(ex_mem_offset[16]), .A3(n194), .A4(
        id_mem_offset[16]), .Y(n98) );
  AO22X1_LVT U71 ( .A1(n189), .A2(ex_mem_offset[15]), .A3(n194), .A4(
        id_mem_offset[15]), .Y(n97) );
  AO22X1_LVT U72 ( .A1(n189), .A2(ex_mem_offset[14]), .A3(n194), .A4(
        id_mem_offset[14]), .Y(n96) );
  AO22X1_LVT U73 ( .A1(n189), .A2(ex_mem_offset[13]), .A3(n194), .A4(
        id_mem_offset[13]), .Y(n95) );
  AO22X1_LVT U74 ( .A1(n189), .A2(ex_mem_offset[12]), .A3(n194), .A4(
        id_mem_offset[12]), .Y(n94) );
  AO22X1_LVT U75 ( .A1(n189), .A2(ex_mem_offset[11]), .A3(n194), .A4(
        id_mem_offset[11]), .Y(n93) );
  AO22X1_LVT U76 ( .A1(n186), .A2(ex_mem_offset[10]), .A3(n191), .A4(
        id_mem_offset[10]), .Y(n92) );
  AO22X1_LVT U77 ( .A1(n186), .A2(ex_mem_offset[9]), .A3(n191), .A4(
        id_mem_offset[9]), .Y(n91) );
  AO22X1_LVT U78 ( .A1(n186), .A2(ex_mem_offset[8]), .A3(n191), .A4(
        id_mem_offset[8]), .Y(n90) );
  AO22X1_LVT U79 ( .A1(n186), .A2(ex_mem_offset[7]), .A3(n191), .A4(
        id_mem_offset[7]), .Y(n89) );
  AO22X1_LVT U80 ( .A1(n186), .A2(ex_mem_offset[6]), .A3(n191), .A4(
        id_mem_offset[6]), .Y(n88) );
  AO22X1_LVT U81 ( .A1(n186), .A2(ex_mem_offset[5]), .A3(n191), .A4(
        id_mem_offset[5]), .Y(n87) );
  AO22X1_LVT U84 ( .A1(n186), .A2(ex_mem_offset[4]), .A3(n191), .A4(
        id_mem_offset[4]), .Y(n86) );
  AO22X1_LVT U85 ( .A1(n186), .A2(ex_mem_offset[3]), .A3(n191), .A4(
        id_mem_offset[3]), .Y(n85) );
  AO22X1_LVT U86 ( .A1(n186), .A2(ex_mem_offset[2]), .A3(n191), .A4(
        id_mem_offset[2]), .Y(n84) );
  AO22X1_LVT U87 ( .A1(n186), .A2(ex_mem_offset[1]), .A3(n191), .A4(
        id_mem_offset[1]), .Y(n83) );
  AO22X1_LVT U88 ( .A1(n186), .A2(ex_mem_offset[0]), .A3(n191), .A4(
        id_mem_offset[0]), .Y(n82) );
  AO22X1_LVT U89 ( .A1(n186), .A2(ex_aluop[4]), .A3(n191), .A4(id_aluop[4]), 
        .Y(n81) );
  AO22X1_LVT U90 ( .A1(n186), .A2(ex_aluop[3]), .A3(n191), .A4(id_aluop[3]), 
        .Y(n80) );
  AO22X1_LVT U91 ( .A1(n186), .A2(ex_aluop[2]), .A3(n191), .A4(id_aluop[2]), 
        .Y(n79) );
  AO22X1_LVT U92 ( .A1(n186), .A2(ex_aluop[1]), .A3(n191), .A4(id_aluop[1]), 
        .Y(n78) );
  AO22X1_LVT U93 ( .A1(n186), .A2(ex_aluop[0]), .A3(n191), .A4(id_aluop[0]), 
        .Y(n77) );
  AO22X1_LVT U94 ( .A1(n186), .A2(ex_alusel[2]), .A3(n191), .A4(id_alusel[2]), 
        .Y(n76) );
  AO22X1_LVT U95 ( .A1(n186), .A2(ex_alusel[1]), .A3(n191), .A4(id_alusel[1]), 
        .Y(n75) );
  AO22X1_LVT U100 ( .A1(n186), .A2(ex_alusel[0]), .A3(n191), .A4(id_alusel[0]), 
        .Y(n74) );
  AO22X1_LVT U101 ( .A1(n186), .A2(ex_opv1[31]), .A3(n191), .A4(id_opv1[31]), 
        .Y(n73) );
  AO22X1_LVT U102 ( .A1(n186), .A2(ex_opv1[30]), .A3(n191), .A4(id_opv1[30]), 
        .Y(n72) );
  AO22X1_LVT U103 ( .A1(n186), .A2(ex_opv1[29]), .A3(n191), .A4(id_opv1[29]), 
        .Y(n71) );
  AO22X1_LVT U104 ( .A1(n186), .A2(ex_opv1[28]), .A3(n191), .A4(id_opv1[28]), 
        .Y(n70) );
  AO22X1_LVT U105 ( .A1(n189), .A2(ex_opv1[27]), .A3(n194), .A4(id_opv1[27]), 
        .Y(n69) );
  AO22X1_LVT U106 ( .A1(n189), .A2(ex_opv1[26]), .A3(n194), .A4(id_opv1[26]), 
        .Y(n68) );
  AO22X1_LVT U107 ( .A1(n189), .A2(ex_opv1[25]), .A3(n194), .A4(id_opv1[25]), 
        .Y(n67) );
  AO22X1_LVT U108 ( .A1(n189), .A2(ex_opv1[24]), .A3(n194), .A4(id_opv1[24]), 
        .Y(n66) );
  AO22X1_LVT U109 ( .A1(n189), .A2(ex_opv1[23]), .A3(n194), .A4(id_opv1[23]), 
        .Y(n65) );
  AO22X1_LVT U110 ( .A1(n189), .A2(ex_opv1[22]), .A3(n194), .A4(id_opv1[22]), 
        .Y(n64) );
  AO22X1_LVT U111 ( .A1(n189), .A2(ex_opv1[21]), .A3(n194), .A4(id_opv1[21]), 
        .Y(n63) );
  AO22X1_LVT U114 ( .A1(n189), .A2(ex_opv1[20]), .A3(n194), .A4(id_opv1[20]), 
        .Y(n62) );
  AO22X1_LVT U115 ( .A1(n189), .A2(ex_opv1[19]), .A3(n194), .A4(id_opv1[19]), 
        .Y(n61) );
  AO22X1_LVT U116 ( .A1(n189), .A2(ex_opv1[18]), .A3(n194), .A4(id_opv1[18]), 
        .Y(n60) );
  AO22X1_LVT U117 ( .A1(n189), .A2(ex_opv1[17]), .A3(n194), .A4(id_opv1[17]), 
        .Y(n59) );
  AO22X1_LVT U118 ( .A1(n189), .A2(ex_opv1[16]), .A3(n194), .A4(id_opv1[16]), 
        .Y(n58) );
  AO22X1_LVT U119 ( .A1(n189), .A2(ex_opv1[15]), .A3(n194), .A4(id_opv1[15]), 
        .Y(n57) );
  AO22X1_LVT U120 ( .A1(n189), .A2(ex_opv1[14]), .A3(n194), .A4(id_opv1[14]), 
        .Y(n56) );
  AO22X1_LVT U121 ( .A1(n190), .A2(ex_opv1[13]), .A3(n195), .A4(id_opv1[13]), 
        .Y(n55) );
  AO22X1_LVT U122 ( .A1(n190), .A2(ex_opv1[12]), .A3(n195), .A4(id_opv1[12]), 
        .Y(n54) );
  AO22X1_LVT U123 ( .A1(n189), .A2(ex_opv1[11]), .A3(n194), .A4(id_opv1[11]), 
        .Y(n53) );
  AO22X1_LVT U124 ( .A1(n189), .A2(ex_opv1[10]), .A3(n194), .A4(id_opv1[10]), 
        .Y(n52) );
  AO22X1_LVT U125 ( .A1(n189), .A2(ex_opv1[9]), .A3(n194), .A4(id_opv1[9]), 
        .Y(n51) );
  AO22X1_LVT U128 ( .A1(n190), .A2(ex_opv1[8]), .A3(n195), .A4(id_opv1[8]), 
        .Y(n50) );
  AO22X1_LVT U129 ( .A1(n190), .A2(ex_opv1[7]), .A3(n195), .A4(id_opv1[7]), 
        .Y(n49) );
  AO22X1_LVT U130 ( .A1(n190), .A2(ex_opv1[6]), .A3(n195), .A4(id_opv1[6]), 
        .Y(n48) );
  AO22X1_LVT U131 ( .A1(n190), .A2(ex_opv1[5]), .A3(n195), .A4(id_opv1[5]), 
        .Y(n47) );
  AO22X1_LVT U132 ( .A1(n186), .A2(ex_opv1[4]), .A3(n191), .A4(id_opv1[4]), 
        .Y(n46) );
  AO22X1_LVT U133 ( .A1(n186), .A2(ex_opv1[3]), .A3(n191), .A4(id_opv1[3]), 
        .Y(n45) );
  AO22X1_LVT U134 ( .A1(n186), .A2(ex_opv1[2]), .A3(n191), .A4(id_opv1[2]), 
        .Y(n44) );
  AO22X1_LVT U135 ( .A1(n186), .A2(ex_opv1[1]), .A3(n191), .A4(id_opv1[1]), 
        .Y(n43) );
  AO22X1_LVT U136 ( .A1(n186), .A2(ex_opv1[0]), .A3(n191), .A4(id_opv1[0]), 
        .Y(n42) );
  AO22X1_LVT U137 ( .A1(n190), .A2(ex_opv2[31]), .A3(n195), .A4(id_opv2[31]), 
        .Y(n41) );
  AO22X1_LVT U138 ( .A1(n190), .A2(ex_opv2[30]), .A3(n195), .A4(id_opv2[30]), 
        .Y(n40) );
  AO22X1_LVT U139 ( .A1(n190), .A2(ex_opv2[29]), .A3(n195), .A4(id_opv2[29]), 
        .Y(n39) );
  AO22X1_LVT U146 ( .A1(n188), .A2(ex_opv2[28]), .A3(n193), .A4(id_opv2[28]), 
        .Y(n38) );
  AO22X1_LVT U147 ( .A1(n188), .A2(ex_opv2[27]), .A3(n193), .A4(id_opv2[27]), 
        .Y(n37) );
  AO22X1_LVT U148 ( .A1(n188), .A2(ex_opv2[26]), .A3(n193), .A4(id_opv2[26]), 
        .Y(n36) );
  AO22X1_LVT U149 ( .A1(n188), .A2(ex_opv2[25]), .A3(n193), .A4(id_opv2[25]), 
        .Y(n35) );
  AO22X1_LVT U150 ( .A1(n188), .A2(ex_opv2[24]), .A3(n193), .A4(id_opv2[24]), 
        .Y(n34) );
  AO22X1_LVT U151 ( .A1(n188), .A2(ex_opv2[23]), .A3(n193), .A4(id_opv2[23]), 
        .Y(n33) );
  AO22X1_LVT U152 ( .A1(n188), .A2(ex_opv2[22]), .A3(n193), .A4(id_opv2[22]), 
        .Y(n32) );
  AO22X1_LVT U153 ( .A1(n188), .A2(ex_opv2[21]), .A3(n193), .A4(id_opv2[21]), 
        .Y(n31) );
  AO22X1_LVT U154 ( .A1(n188), .A2(ex_opv2[20]), .A3(n193), .A4(id_opv2[20]), 
        .Y(n30) );
  AO22X1_LVT U155 ( .A1(n188), .A2(ex_opv2[19]), .A3(n193), .A4(id_opv2[19]), 
        .Y(n29) );
  AO22X1_LVT U156 ( .A1(n188), .A2(ex_opv2[18]), .A3(n193), .A4(id_opv2[18]), 
        .Y(n28) );
  AO22X1_LVT U157 ( .A1(n188), .A2(ex_opv2[17]), .A3(n193), .A4(id_opv2[17]), 
        .Y(n27) );
  AO22X1_LVT U160 ( .A1(n188), .A2(ex_opv2[16]), .A3(n193), .A4(id_opv2[16]), 
        .Y(n26) );
  AO22X1_LVT U161 ( .A1(n188), .A2(ex_opv2[15]), .A3(n193), .A4(id_opv2[15]), 
        .Y(n25) );
  AO22X1_LVT U162 ( .A1(n188), .A2(ex_opv2[14]), .A3(n193), .A4(id_opv2[14]), 
        .Y(n24) );
  AO22X1_LVT U163 ( .A1(n188), .A2(ex_opv2[13]), .A3(n193), .A4(id_opv2[13]), 
        .Y(n23) );
  AO22X1_LVT U164 ( .A1(n188), .A2(ex_opv2[12]), .A3(n193), .A4(id_opv2[12]), 
        .Y(n22) );
  AO22X1_LVT U165 ( .A1(n188), .A2(ex_opv2[11]), .A3(n193), .A4(id_opv2[11]), 
        .Y(n21) );
  AO22X1_LVT U166 ( .A1(n188), .A2(ex_opv2[10]), .A3(n193), .A4(id_opv2[10]), 
        .Y(n20) );
  AO22X1_LVT U167 ( .A1(n188), .A2(ex_opv2[9]), .A3(n193), .A4(id_opv2[9]), 
        .Y(n19) );
  AO22X1_LVT U168 ( .A1(n188), .A2(ex_opv2[8]), .A3(n193), .A4(id_opv2[8]), 
        .Y(n18) );
  AO22X1_LVT U169 ( .A1(n188), .A2(ex_opv2[7]), .A3(n193), .A4(id_opv2[7]), 
        .Y(n17) );
  AO22X1_LVT U170 ( .A1(n188), .A2(ex_opv2[6]), .A3(n193), .A4(id_opv2[6]), 
        .Y(n16) );
  AO22X1_LVT U171 ( .A1(n188), .A2(ex_opv2[5]), .A3(n193), .A4(id_opv2[5]), 
        .Y(n15) );
  AO22X1_LVT U174 ( .A1(n190), .A2(ex_opv2[4]), .A3(n195), .A4(id_opv2[4]), 
        .Y(n14) );
  AO22X1_LVT U175 ( .A1(n190), .A2(ex_opv2[3]), .A3(n195), .A4(id_opv2[3]), 
        .Y(n13) );
  AO22X1_LVT U176 ( .A1(n190), .A2(ex_opv2[2]), .A3(n195), .A4(id_opv2[2]), 
        .Y(n12) );
  AO22X1_LVT U177 ( .A1(n190), .A2(ex_opv2[1]), .A3(n195), .A4(id_opv2[1]), 
        .Y(n11) );
  AO22X1_LVT U178 ( .A1(n190), .A2(ex_opv2[0]), .A3(n195), .A4(id_opv2[0]), 
        .Y(n10) );
  AO22X1_LVT U179 ( .A1(n186), .A2(ex_reg_waddr[4]), .A3(n191), .A4(
        id_reg_waddr[4]), .Y(n9) );
  AO22X1_LVT U180 ( .A1(n186), .A2(ex_reg_waddr[3]), .A3(n191), .A4(
        id_reg_waddr[3]), .Y(n8) );
  AO22X1_LVT U181 ( .A1(n186), .A2(ex_reg_waddr[2]), .A3(n191), .A4(
        id_reg_waddr[2]), .Y(n7) );
  AO22X1_LVT U182 ( .A1(n186), .A2(ex_reg_waddr[1]), .A3(n191), .A4(
        id_reg_waddr[1]), .Y(n6) );
  AO22X1_LVT U183 ( .A1(n186), .A2(ex_reg_waddr[0]), .A3(n191), .A4(
        id_reg_waddr[0]), .Y(n5) );
  INVX1_LVT U3 ( .A(rst), .Y(n185) );
  NBUFFX4_LVT U5 ( .A(n173), .Y(n186) );
  NBUFFX8_LVT U6 ( .A(n173), .Y(n187) );
  NBUFFX4_LVT U7 ( .A(n173), .Y(n188) );
  NBUFFX4_LVT U9 ( .A(n173), .Y(n189) );
  NBUFFX4_LVT U10 ( .A(n173), .Y(n190) );
  NBUFFX4_LVT U11 ( .A(n175), .Y(n191) );
  NBUFFX8_LVT U24 ( .A(n175), .Y(n192) );
  NBUFFX4_LVT U25 ( .A(n175), .Y(n193) );
  NBUFFX4_LVT U38 ( .A(n175), .Y(n194) );
  NBUFFX4_LVT U39 ( .A(n175), .Y(n195) );
  DFFX2_LVT \ex_opv1_reg[3]  ( .D(n45), .CLK(clk), .Q(ex_opv1[3]) );
  DFFX2_LVT \ex_opv1_reg[27]  ( .D(n69), .CLK(clk), .Q(ex_opv1[27]) );
  DFFX2_LVT \ex_opv1_reg[28]  ( .D(n70), .CLK(clk), .Q(ex_opv1[28]) );
  DFFX2_LVT \ex_opv1_reg[5]  ( .D(n47), .CLK(clk), .Q(ex_opv1[5]) );
  DFFX2_LVT \ex_opv1_reg[10]  ( .D(n52), .CLK(clk), .Q(ex_opv1[10]) );
  DFFX2_LVT \ex_opv1_reg[19]  ( .D(n61), .CLK(clk), .Q(ex_opv1[19]) );
  DFFX2_LVT \ex_opv1_reg[13]  ( .D(n55), .CLK(clk), .Q(ex_opv1[13]) );
  DFFX2_LVT \ex_opv1_reg[17]  ( .D(n59), .CLK(clk), .Q(ex_opv1[17]) );
  DFFX2_LVT \ex_opv1_reg[11]  ( .D(n53), .CLK(clk), .Q(ex_opv1[11]) );
  DFFX2_LVT \ex_opv1_reg[26]  ( .D(n68), .CLK(clk), .Q(ex_opv1[26]) );
  DFFX2_LVT \ex_opv1_reg[30]  ( .D(n72), .CLK(clk), .Q(ex_opv1[30]) );
  DFFX2_LVT \ex_opv1_reg[18]  ( .D(n60), .CLK(clk), .Q(ex_opv1[18]) );
  DFFX2_LVT \ex_opv1_reg[20]  ( .D(n62), .CLK(clk), .Q(ex_opv1[20]) );
  DFFX2_LVT \ex_opv1_reg[9]  ( .D(n51), .CLK(clk), .Q(ex_opv1[9]) );
  DFFX2_LVT \ex_opv1_reg[8]  ( .D(n50), .CLK(clk), .Q(ex_opv1[8]) );
  DFFX2_LVT \ex_opv1_reg[16]  ( .D(n58), .CLK(clk), .Q(ex_opv1[16]) );
  DFFX2_LVT \ex_opv1_reg[7]  ( .D(n49), .CLK(clk), .Q(ex_opv1[7]) );
  DFFX2_LVT \ex_opv1_reg[2]  ( .D(n44), .CLK(clk), .Q(ex_opv1[2]) );
  DFFX2_LVT \ex_opv1_reg[6]  ( .D(n48), .CLK(clk), .Q(ex_opv1[6]) );
  DFFX2_LVT \ex_opv1_reg[4]  ( .D(n46), .CLK(clk), .Q(ex_opv1[4]) );
  DFFX2_LVT \ex_opv1_reg[25]  ( .D(n67), .CLK(clk), .Q(ex_opv1[25]) );
  DFFX2_LVT \ex_opv2_reg[9]  ( .D(n19), .CLK(clk), .Q(ex_opv2[9]) );
  DFFX2_LVT \ex_aluop_reg[1]  ( .D(n78), .CLK(clk), .Q(ex_aluop[1]) );
  DFFX2_LVT \ex_aluop_reg[2]  ( .D(n79), .CLK(clk), .Q(ex_aluop[2]) );
  DFFX2_LVT \ex_aluop_reg[4]  ( .D(n81), .CLK(clk), .Q(ex_aluop[4]) );
  DFFX2_LVT ex_we_reg ( .D(n146), .CLK(clk), .Q(ex_we) );
  DFFX1_LVT \ex_opv1_reg[29]  ( .D(n71), .CLK(clk), .Q(ex_opv1[29]) );
  DFFX1_LVT \ex_opv1_reg[31]  ( .D(n73), .CLK(clk), .Q(ex_opv1[31]) );
  DFFX1_LVT \ex_opv1_reg[15]  ( .D(n57), .CLK(clk), .Q(ex_opv1[15]) );
  DFFX1_LVT \ex_opv1_reg[14]  ( .D(n56), .CLK(clk), .Q(ex_opv1[14]) );
  DFFX1_LVT \ex_opv1_reg[21]  ( .D(n63), .CLK(clk), .Q(ex_opv1[21]) );
  DFFX1_LVT \ex_opv1_reg[24]  ( .D(n66), .CLK(clk), .Q(ex_opv1[24]) );
  DFFX1_LVT \ex_opv1_reg[12]  ( .D(n54), .CLK(clk), .Q(ex_opv1[12]) );
  DFFX1_LVT \ex_opv1_reg[22]  ( .D(n64), .CLK(clk), .Q(ex_opv1[22]) );
  DFFX1_LVT \ex_opv1_reg[1]  ( .D(n43), .CLK(clk), .Q(ex_opv1[1]) );
  DFFX1_LVT \ex_opv1_reg[23]  ( .D(n65), .CLK(clk), .Q(ex_opv1[23]) );
endmodule


module execute_alu ( rst, aluop, alusel, opv1, opv2, reg_waddr_i, we_i, 
        link_addr, mem_offset, reg_waddr_o, we_o, reg_wdata, stallreq, 
        mem_addr, ex_aluop, rt_data );
  input [7:0] aluop;
  input [2:0] alusel;
  input [31:0] opv1;
  input [31:0] opv2;
  input [4:0] reg_waddr_i;
  input [31:0] link_addr;
  input [31:0] mem_offset;
  output [4:0] reg_waddr_o;
  output [31:0] reg_wdata;
  output [31:0] mem_addr;
  output [7:0] ex_aluop;
  output [31:0] rt_data;
  input rst, we_i;
  output we_o, stallreq;
  wire   we_i, N287, n2, n4, n5, n6, n8, n10, n13, n14, n15, n16, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n37, n38, n41, n42, n43, n44, n45, n46, n48, n49, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n76, n77, n81, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n97, n98, n100, n101, n104, n105,
         n106, n107, n108, n109, n111, n113, n115, n116, n117, n119, n120,
         n121, n122, n123, n125, n126, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n150, n151, n152, n153, n154, n155, n156, n157, n160,
         n161, n162, n163, n166, n167, n168, n169, n172, n173, n174, n175,
         n176, n177, n178, n179, n181, n182, n184, n185, n188, n190, n192,
         n194, n195, n196, n197, n198, n199, n200, n202, n203, n204, n205,
         n206, n207, n208, n209, n211, n212, n215, n216, n217, n218, n219,
         n221, n222, n223, n224, n225, n226, n227, n229, n230, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n244, n245, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n270, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n284,
         n285, n286, n288, n289, n291, n292, n293, n294, n295, n296, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n334, n335, n336,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n358, n359, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n430,
         n431, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n507, n508, n509, n510, n511,
         n513, n514, n515, n516, n517, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n562, n563, n564, n565, n568, n569, n570, n571, n573, n574,
         n575, n576, n577, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n594, n596, n597, n598, n599, n600,
         n601, n602, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n667, n668, n669, n671,
         n672, n673, n674, n675, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n753, n754, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n769, n770, n771, n772, n773, n774, n776, n777, n778, n779, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n829,
         n830, n831, n833, n834, n836, n837, n838, n839, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n875, n876, n877, n878, n879,
         n880, n881, n883, n884, n885, n886, n887, n888, n890, n891, n892,
         n893, n894, n895, n896, n897, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n919, n920, n921, n925, n926, n927, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n939, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n968,
         n969, n970, n971, n972, n973, n975, n976, n977, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n991, n992, n993,
         n994, n996, n998, n999, n1001, n1002, n1004, n1005, n1006, n1007,
         n1009, n1010, n1011, n1012, n1013, n1014, n1016, n1018, n1019, n1020,
         n1021, n1023, n1026, n1028, n1030, n1031, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1139, n1140, n1141, n1142, n1143, n1144;
  assign reg_waddr_o[4] = reg_waddr_i[4];
  assign reg_waddr_o[3] = reg_waddr_i[3];
  assign reg_waddr_o[2] = reg_waddr_i[2];
  assign reg_waddr_o[1] = reg_waddr_i[1];
  assign reg_waddr_o[0] = reg_waddr_i[0];
  assign we_o = we_i;
  assign ex_aluop[4] = aluop[4];
  assign ex_aluop[3] = aluop[3];
  assign ex_aluop[2] = aluop[2];
  assign ex_aluop[1] = aluop[1];
  assign rt_data[31] = opv2[31];
  assign rt_data[30] = opv2[30];
  assign rt_data[29] = opv2[29];
  assign rt_data[28] = opv2[28];
  assign rt_data[27] = opv2[27];
  assign rt_data[26] = opv2[26];
  assign rt_data[25] = opv2[25];
  assign rt_data[24] = opv2[24];
  assign rt_data[23] = opv2[23];
  assign rt_data[22] = opv2[22];
  assign rt_data[21] = opv2[21];
  assign rt_data[20] = opv2[20];
  assign rt_data[19] = opv2[19];
  assign rt_data[18] = opv2[18];
  assign rt_data[17] = opv2[17];
  assign rt_data[16] = opv2[16];
  assign rt_data[15] = opv2[15];
  assign rt_data[14] = opv2[14];
  assign rt_data[13] = opv2[13];
  assign rt_data[12] = opv2[12];
  assign rt_data[11] = opv2[11];
  assign rt_data[10] = opv2[10];
  assign rt_data[8] = opv2[8];
  assign rt_data[7] = opv2[7];
  assign rt_data[6] = opv2[6];
  assign rt_data[5] = opv2[5];
  assign rt_data[4] = opv2[4];
  assign rt_data[3] = opv2[3];
  assign rt_data[2] = opv2[2];
  assign rt_data[1] = opv2[1];
  assign rt_data[0] = N287;
  assign N287 = opv2[0];

  NOR4X1_LVT U6 ( .A1(aluop[2]), .A2(rst), .A3(aluop[4]), .A4(alusel[1]), .Y(
        n37) );
  INVX1_LVT U7 ( .A(alusel[0]), .Y(n48) );
  AND4X1_LVT U8 ( .A1(aluop[3]), .A2(alusel[2]), .A3(n37), .A4(n48), .Y(n248)
         );
  INVX1_LVT U9 ( .A(n248), .Y(n6) );
  NOR2X0_LVT U14 ( .A1(n1031), .A2(aluop[1]), .Y(n4) );
  NOR2X0_LVT U15 ( .A1(n1139), .A2(n4), .Y(n5) );
  XOR2X1_LVT U19 ( .A1(n1139), .A2(opv2[30]), .Y(n560) );
  XOR2X1_LVT U20 ( .A1(n1139), .A2(opv2[29]), .Y(n989) );
  XOR2X1_LVT U21 ( .A1(n1139), .A2(opv2[28]), .Y(n527) );
  XOR2X1_LVT U22 ( .A1(n1139), .A2(opv2[27]), .Y(n959) );
  XOR2X1_LVT U23 ( .A1(n1139), .A2(opv2[26]), .Y(n936) );
  XOR2X1_LVT U24 ( .A1(n1139), .A2(opv2[25]), .Y(n489) );
  XOR2X1_LVT U25 ( .A1(n1139), .A2(opv2[24]), .Y(n444) );
  XOR2X1_LVT U26 ( .A1(n1139), .A2(opv2[23]), .Y(n407) );
  XOR2X1_LVT U27 ( .A1(n1139), .A2(opv2[22]), .Y(n384) );
  XOR2X1_LVT U28 ( .A1(n1139), .A2(opv2[21]), .Y(n908) );
  XOR2X1_LVT U29 ( .A1(n1139), .A2(opv2[20]), .Y(n885) );
  XOR2X1_LVT U30 ( .A1(n1139), .A2(opv2[19]), .Y(n865) );
  XOR2X1_LVT U31 ( .A1(n1139), .A2(opv2[18]), .Y(n369) );
  XOR2X1_LVT U32 ( .A1(n1139), .A2(opv2[17]), .Y(n845) );
  XOR2X1_LVT U33 ( .A1(n1139), .A2(opv2[16]), .Y(n819) );
  XOR2X1_LVT U34 ( .A1(n1139), .A2(opv2[15]), .Y(n791) );
  XOR2X1_LVT U35 ( .A1(n1139), .A2(opv2[14]), .Y(n345) );
  XOR2X1_LVT U36 ( .A1(n1139), .A2(opv2[13]), .Y(n767) );
  XOR2X1_LVT U37 ( .A1(n2), .A2(opv2[12]), .Y(n745) );
  XOR2X1_LVT U38 ( .A1(n2), .A2(opv2[11]), .Y(n729) );
  XOR2X1_LVT U39 ( .A1(n2), .A2(opv2[10]), .Y(n54) );
  XOR2X1_LVT U40 ( .A1(n2), .A2(opv2[9]), .Y(n92) );
  XOR2X1_LVT U41 ( .A1(n2), .A2(opv2[8]), .Y(n711) );
  XOR2X1_LVT U42 ( .A1(n2), .A2(opv2[7]), .Y(n116) );
  XOR2X1_LVT U44 ( .A1(n2), .A2(opv2[6]), .Y(n326) );
  XOR2X1_LVT U45 ( .A1(n2), .A2(opv2[5]), .Y(n693) );
  XOR2X1_LVT U46 ( .A1(n2), .A2(opv2[4]), .Y(n675) );
  XOR2X1_LVT U47 ( .A1(n2), .A2(opv2[3]), .Y(n305) );
  XOR2X1_LVT U48 ( .A1(n2), .A2(opv2[2]), .Y(n280) );
  XOR2X1_LVT U49 ( .A1(n2), .A2(opv2[1]), .Y(n254) );
  XOR2X1_LVT U50 ( .A1(n2), .A2(N287), .Y(n133) );
  NOR4X1_LVT U51 ( .A1(aluop[3]), .A2(alusel[2]), .A3(rst), .A4(aluop[4]), .Y(
        n8) );
  NAND2X0_LVT U56 ( .A1(n1035), .A2(n1036), .Y(n176) );
  NAND3X0_LVT U62 ( .A1(n1085), .A2(n1040), .A3(n1038), .Y(n88) );
  NAND2X0_LVT U65 ( .A1(n1001), .A2(n1042), .Y(n587) );
  INVX1_LVT U66 ( .A(n587), .Y(n10) );
  NOR3X0_LVT U67 ( .A1(n1081), .A2(n1089), .A3(n10), .Y(n987) );
  NAND2X0_LVT U70 ( .A1(aluop[1]), .A2(n430), .Y(n588) );
  INVX1_LVT U71 ( .A(n588), .Y(n350) );
  NAND2X0_LVT U72 ( .A1(n350), .A2(n1042), .Y(n812) );
  NAND2X0_LVT U74 ( .A1(n28), .A2(n1090), .Y(n807) );
  INVX2_LVT U75 ( .A(n807), .Y(n985) );
  AO22X1_LVT U76 ( .A1(N287), .A2(n1143), .A3(n1035), .A4(opv1[30]), .Y(n139)
         );
  AND2X1_LVT U77 ( .A1(n1036), .A2(n139), .Y(n351) );
  AND2X1_LVT U81 ( .A1(opv2[2]), .A2(n1040), .Y(n13) );
  NAND2X0_LVT U86 ( .A1(opv1[25]), .A2(n16), .Y(n141) );
  NAND2X0_LVT U87 ( .A1(N287), .A2(opv2[1]), .Y(n86) );
  NAND2X0_LVT U90 ( .A1(n1112), .A2(n1080), .Y(n135) );
  NAND2X0_LVT U91 ( .A1(n1085), .A2(opv1[26]), .Y(n14) );
  NAND2X0_LVT U92 ( .A1(opv2[1]), .A2(n1035), .Y(n29) );
  NAND2X0_LVT U95 ( .A1(n1115), .A2(n1082), .Y(n62) );
  NAND4X0_LVT U96 ( .A1(n141), .A2(n135), .A3(n14), .A4(n62), .Y(n934) );
  NAND2X0_LVT U101 ( .A1(n1119), .A2(n16), .Y(n136) );
  NAND2X0_LVT U103 ( .A1(n1135), .A2(n1080), .Y(n137) );
  NAND2X0_LVT U105 ( .A1(n1085), .A2(n1113), .Y(n63) );
  NAND2X0_LVT U106 ( .A1(n1128), .A2(n1082), .Y(n59) );
  NAND4X0_LVT U107 ( .A1(n136), .A2(n137), .A3(n63), .A4(n59), .Y(n947) );
  AO22X1_LVT U108 ( .A1(n1084), .A2(n934), .A3(n15), .A4(n947), .Y(n18) );
  INVX1_LVT U109 ( .A(n18), .Y(n26) );
  NAND2X0_LVT U113 ( .A1(n1133), .A2(n16), .Y(n138) );
  NAND2X0_LVT U114 ( .A1(n1120), .A2(n1080), .Y(n143) );
  NAND2X0_LVT U115 ( .A1(n1085), .A2(n1130), .Y(n60) );
  NAND2X0_LVT U116 ( .A1(n1127), .A2(n1082), .Y(n57) );
  NAND4X0_LVT U117 ( .A1(n138), .A2(n143), .A3(n60), .A4(n57), .Y(n946) );
  AO22X1_LVT U118 ( .A1(n1001), .A2(n1131), .A3(n19), .A4(n946), .Y(n20) );
  INVX1_LVT U119 ( .A(n20), .Y(n25) );
  NAND2X0_LVT U120 ( .A1(opv1[29]), .A2(n16), .Y(n22) );
  NAND2X0_LVT U121 ( .A1(n1080), .A2(opv1[27]), .Y(n142) );
  NAND2X0_LVT U122 ( .A1(n1140), .A2(n1082), .Y(n21) );
  NAND3X0_LVT U123 ( .A1(n22), .A2(n142), .A3(n21), .Y(n23) );
  NAND2X0_LVT U124 ( .A1(n28), .A2(n23), .Y(n24) );
  NAND3X0_LVT U125 ( .A1(n26), .A2(n25), .A3(n24), .Y(n31) );
  NAND2X0_LVT U127 ( .A1(n1031), .A2(n1034), .Y(n389) );
  INVX1_LVT U128 ( .A(n389), .Y(n27) );
  NAND3X0_LVT U129 ( .A1(n27), .A2(n430), .A3(opv2[4]), .Y(n976) );
  INVX2_LVT U130 ( .A(n976), .Y(n1013) );
  NAND2X0_LVT U131 ( .A1(n1080), .A2(n1126), .Y(n147) );
  NAND2X0_LVT U132 ( .A1(n1123), .A2(n16), .Y(n146) );
  NAND2X0_LVT U133 ( .A1(n1129), .A2(n1082), .Y(n288) );
  NAND2X0_LVT U134 ( .A1(n1085), .A2(n1136), .Y(n56) );
  NAND4X0_LVT U135 ( .A1(n147), .A2(n146), .A3(n288), .A4(n56), .Y(n387) );
  NAND2X0_LVT U137 ( .A1(n1134), .A2(n16), .Y(n144) );
  NAND2X0_LVT U138 ( .A1(n1132), .A2(n1080), .Y(n145) );
  NAND2X0_LVT U139 ( .A1(n1085), .A2(n1117), .Y(n58) );
  NAND2X0_LVT U140 ( .A1(n1116), .A2(n1082), .Y(n55) );
  NAND4X0_LVT U141 ( .A1(n144), .A2(n145), .A3(n58), .A4(n55), .Y(n945) );
  OA22X1_LVT U145 ( .A1(n1037), .A2(n29), .A3(n176), .A4(n1041), .Y(n30) );
  NAND2X0_LVT U146 ( .A1(opv1[1]), .A2(n16), .Y(n151) );
  NAND2X0_LVT U147 ( .A1(n30), .A2(n151), .Y(n373) );
  NAND2X0_LVT U148 ( .A1(n1137), .A2(n16), .Y(n148) );
  NAND2X0_LVT U149 ( .A1(n1142), .A2(n1080), .Y(n150) );
  NAND2X0_LVT U150 ( .A1(n1085), .A2(n1125), .Y(n289) );
  NAND2X0_LVT U151 ( .A1(n1114), .A2(n1082), .Y(n291) );
  NAND4X0_LVT U152 ( .A1(n148), .A2(n150), .A3(n289), .A4(n291), .Y(n374) );
  AO22X1_LVT U153 ( .A1(opv2[2]), .A2(n373), .A3(n1038), .A4(n374), .Y(n386)
         );
  AO222X1_LVT U154 ( .A1(n387), .A2(n1084), .A3(n945), .A4(n28), .A5(n386), 
        .A6(opv2[3]), .Y(n358) );
  AO22X1_LVT U155 ( .A1(n1086), .A2(n31), .A3(n1013), .A4(n358), .Y(n32) );
  AO21X1_LVT U156 ( .A1(n985), .A2(n351), .A3(n32), .Y(n33) );
  AO21X1_LVT U157 ( .A1(n987), .A2(n1143), .A3(n33), .Y(n34) );
  INVX1_LVT U160 ( .A(n37), .Y(n38) );
  NOR4X1_LVT U161 ( .A1(n48), .A2(n38), .A3(alusel[2]), .A4(aluop[3]), .Y(n65)
         );
  OR2X1_LVT U167 ( .A1(n1078), .A2(n1131), .Y(n234) );
  INVX1_LVT U168 ( .A(n234), .Y(n46) );
  AND2X1_LVT U169 ( .A1(n1131), .A2(n1078), .Y(n230) );
  AND2X1_LVT U170 ( .A1(opv2[30]), .A2(n1131), .Y(n44) );
  NAND2X0_LVT U171 ( .A1(n1088), .A2(n1033), .Y(n972) );
  INVX1_LVT U172 ( .A(n972), .Y(n529) );
  INVX1_LVT U173 ( .A(n529), .Y(n42) );
  NAND3X0_LVT U174 ( .A1(ex_aluop[0]), .A2(n65), .A3(n1034), .Y(n973) );
  INVX1_LVT U175 ( .A(n973), .Y(n546) );
  INVX1_LVT U176 ( .A(n546), .Y(n41) );
  NAND2X0_LVT U177 ( .A1(n42), .A2(n41), .Y(n43) );
  AND2X1_LVT U178 ( .A1(n44), .A2(n43), .Y(n45) );
  NAND2X0_LVT U183 ( .A1(n66), .A2(link_addr[30]), .Y(n49) );
  NAND3X0_LVT U184 ( .A1(n1111), .A2(n1110), .A3(n49), .Y(reg_wdata[30]) );
  FADDX1_LVT U186 ( .A(opv1[10]), .B(n54), .CI(n53), .CO(n728), .S(n74) );
  NAND2X0_LVT U187 ( .A1(n1134), .A2(n1080), .Y(n467) );
  NAND2X0_LVT U188 ( .A1(n1132), .A2(n16), .Y(n471) );
  NAND4X0_LVT U189 ( .A1(n56), .A2(n55), .A3(n467), .A4(n471), .Y(n334) );
  NAND2X0_LVT U190 ( .A1(n985), .A2(n334), .Y(n72) );
  AOI222X1_LVT U192 ( .A1(n374), .A2(n1084), .A3(n387), .A4(n28), .A5(n373), 
        .A6(n15), .Y(n949) );
  NAND2X0_LVT U193 ( .A1(n1120), .A2(n16), .Y(n468) );
  NAND2X0_LVT U194 ( .A1(n1133), .A2(n1080), .Y(n475) );
  NAND4X0_LVT U195 ( .A1(n58), .A2(n57), .A3(n468), .A4(n475), .Y(n346) );
  NAND2X0_LVT U196 ( .A1(n1135), .A2(n16), .Y(n476) );
  NAND2X0_LVT U197 ( .A1(n1119), .A2(n1080), .Y(n448) );
  NAND4X0_LVT U198 ( .A1(n60), .A2(n59), .A3(n476), .A4(n448), .Y(n347) );
  NAND2X0_LVT U200 ( .A1(n1080), .A2(n1121), .Y(n537) );
  NAND2X0_LVT U201 ( .A1(n1112), .A2(n16), .Y(n449) );
  NAND4X0_LVT U202 ( .A1(n63), .A2(n62), .A3(n537), .A4(n449), .Y(n349) );
  AOI222X1_LVT U203 ( .A1(n346), .A2(n1083), .A3(n347), .A4(n15), .A5(n349), 
        .A6(n19), .Y(n64) );
  OA22X1_LVT U204 ( .A1(n949), .A2(n1118), .A3(n64), .A4(n812), .Y(n71) );
  NAND2X0_LVT U205 ( .A1(n65), .A2(n1034), .Y(n798) );
  NAND4X0_LVT U207 ( .A1(n1031), .A2(n1136), .A3(opv2[10]), .A4(n1087), .Y(n70) );
  NAND3X0_LVT U210 ( .A1(n1031), .A2(n1136), .A3(opv2[10]), .Y(n67) );
  OA21X1_LVT U211 ( .A1(n1136), .A2(opv2[10]), .A3(n67), .Y(n68) );
  AOI22X1_LVT U212 ( .A1(n66), .A2(link_addr[10]), .A3(n1088), .A4(n68), .Y(
        n69) );
  NAND4X0_LVT U213 ( .A1(n72), .A2(n71), .A3(n70), .A4(n69), .Y(n73) );
  AND4X1_LVT U216 ( .A1(n430), .A2(opv2[4]), .A3(n1139), .A4(n88), .Y(n777) );
  OA221X1_LVT U217 ( .A1(n1085), .A2(opv2[2]), .A3(n176), .A4(n1038), .A5(
        n1143), .Y(n950) );
  NAND2X0_LVT U218 ( .A1(n1085), .A2(n1038), .Y(n464) );
  NAND2X0_LVT U219 ( .A1(opv2[3]), .A2(n464), .Y(n393) );
  NAND2X0_LVT U220 ( .A1(n88), .A2(n393), .Y(n904) );
  AND3X1_LVT U221 ( .A1(n1143), .A2(n777), .A3(n904), .Y(n776) );
  AO21X1_LVT U222 ( .A1(n777), .A2(n950), .A3(n776), .Y(n737) );
  INVX1_LVT U223 ( .A(n737), .Y(n77) );
  MUX41X1_LVT U224 ( .A1(opv1[27]), .A3(n1124), .A2(opv1[29]), .A4(opv1[28]), 
        .S0(n1035), .S1(opv2[1]), .Y(n348) );
  AO22X1_LVT U225 ( .A1(opv2[2]), .A2(n351), .A3(n1038), .A4(n348), .Y(n933)
         );
  AND3X1_LVT U226 ( .A1(opv2[4]), .A2(n350), .A3(n1040), .Y(n732) );
  NAND2X0_LVT U227 ( .A1(n933), .A2(n732), .Y(n76) );
  AOI22X1_LVT U230 ( .A1(n1085), .A2(opv1[29]), .A3(n1143), .A4(n1082), .Y(n81) );
  NAND2X0_LVT U231 ( .A1(opv1[30]), .A2(n16), .Y(n575) );
  NAND2X0_LVT U232 ( .A1(n81), .A2(n575), .Y(n984) );
  NAND2X0_LVT U233 ( .A1(n1124), .A2(n16), .Y(n571) );
  NAND2X0_LVT U234 ( .A1(n1080), .A2(n1140), .Y(n574) );
  NAND2X0_LVT U236 ( .A1(n1141), .A2(n1082), .Y(n1006) );
  NAND2X0_LVT U237 ( .A1(n1085), .A2(n1121), .Y(n516) );
  NAND4X0_LVT U238 ( .A1(n571), .A2(n574), .A3(n1006), .A4(n516), .Y(n784) );
  AO22X1_LVT U239 ( .A1(opv2[2]), .A2(n984), .A3(n1038), .A4(n784), .Y(n520)
         );
  NAND2X0_LVT U240 ( .A1(n1130), .A2(n16), .Y(n425) );
  NAND2X0_LVT U241 ( .A1(n1128), .A2(n1080), .Y(n412) );
  NAND2X0_LVT U242 ( .A1(n1085), .A2(n1133), .Y(n494) );
  NAND2X0_LVT U243 ( .A1(n1135), .A2(n1082), .Y(n502) );
  NAND4X0_LVT U244 ( .A1(n425), .A2(n412), .A3(n494), .A4(n502), .Y(n783) );
  NAND2X0_LVT U245 ( .A1(n1113), .A2(n16), .Y(n413) );
  NAND2X0_LVT U246 ( .A1(n1115), .A2(n1080), .Y(n570) );
  NAND2X0_LVT U247 ( .A1(n1085), .A2(n1119), .Y(n503) );
  NAND2X0_LVT U248 ( .A1(n1112), .A2(n1082), .Y(n515) );
  NAND4X0_LVT U249 ( .A1(n413), .A2(n570), .A3(n503), .A4(n515), .Y(n785) );
  NAND2X0_LVT U251 ( .A1(n1127), .A2(n1080), .Y(n426) );
  NAND2X0_LVT U252 ( .A1(n1117), .A2(n16), .Y(n418) );
  NAND2X0_LVT U253 ( .A1(n1085), .A2(n1134), .Y(n499) );
  NAND2X0_LVT U254 ( .A1(n1120), .A2(n1082), .Y(n495) );
  NAND4X0_LVT U255 ( .A1(n426), .A2(n418), .A3(n499), .A4(n495), .Y(n765) );
  AO222X1_LVT U257 ( .A1(n783), .A2(n15), .A3(n785), .A4(n19), .A5(n765), .A6(
        n1084), .Y(n84) );
  OA222X1_LVT U258 ( .A1(n1042), .A2(n520), .A3(n1042), .A4(n1040), .A5(
        opv2[4]), .A6(n84), .Y(n85) );
  AND2X1_LVT U259 ( .A1(n28), .A2(n1042), .Y(n311) );
  NAND2X0_LVT U260 ( .A1(n1085), .A2(n1123), .Y(n100) );
  NAND2X0_LVT U261 ( .A1(n1136), .A2(n16), .Y(n422) );
  NAND2X0_LVT U262 ( .A1(n1116), .A2(n1080), .Y(n417) );
  NAND2X0_LVT U263 ( .A1(n1132), .A2(n1082), .Y(n498) );
  NAND4X0_LVT U264 ( .A1(n100), .A2(n422), .A3(n417), .A4(n498), .Y(n701) );
  OA221X1_LVT U265 ( .A1(n85), .A2(n311), .A3(n85), .A4(n701), .A5(aluop[1]), 
        .Y(n90) );
  NAND2X0_LVT U266 ( .A1(n176), .A2(n86), .Y(n847) );
  NAND2X0_LVT U267 ( .A1(n950), .A2(n847), .Y(n509) );
  NAND2X0_LVT U268 ( .A1(n1143), .A2(n904), .Y(n87) );
  NAND2X0_LVT U269 ( .A1(n509), .A2(n87), .Y(n708) );
  AND4X1_LVT U270 ( .A1(n1139), .A2(n708), .A3(opv2[4]), .A4(n88), .Y(n89) );
  OR2X1_LVT U271 ( .A1(n90), .A2(n89), .Y(n95) );
  FADDX1_LVT U272 ( .A(opv1[9]), .B(n92), .CI(n91), .CO(n53), .S(n94) );
  NAND3X0_LVT U273 ( .A1(ex_aluop[0]), .A2(n1123), .A3(opv2[9]), .Y(n97) );
  INVX1_LVT U274 ( .A(n97), .Y(n93) );
  OA21X1_LVT U277 ( .A1(n1123), .A2(opv2[9]), .A3(n97), .Y(n98) );
  NAND2X0_LVT U280 ( .A1(n1080), .A2(n1125), .Y(n309) );
  NAND2X0_LVT U281 ( .A1(n1126), .A2(n1082), .Y(n257) );
  NAND2X0_LVT U282 ( .A1(n1129), .A2(n16), .Y(n104) );
  NAND4X0_LVT U283 ( .A1(n309), .A2(n257), .A3(n104), .A4(n100), .Y(n926) );
  AO22X1_LVT U284 ( .A1(opv1[0]), .A2(n16), .A3(n1085), .A4(opv1[1]), .Y(n846)
         );
  MUX41X1_LVT U285 ( .A1(n1114), .A3(n1137), .A2(n1122), .A4(n1142), .S0(n1035), .S1(opv2[1]), .Y(n839) );
  AO222X1_LVT U286 ( .A1(n926), .A2(n28), .A3(n846), .A4(n15), .A5(n839), .A6(
        n1083), .Y(n504) );
  NAND2X0_LVT U287 ( .A1(n1086), .A2(n504), .Y(n101) );
  NAND3X0_LVT U289 ( .A1(n1031), .A2(n1126), .A3(opv2[7]), .Y(n107) );
  INVX1_LVT U290 ( .A(n107), .Y(n105) );
  NAND2X0_LVT U291 ( .A1(n1085), .A2(n1126), .Y(n119) );
  NAND2X0_LVT U292 ( .A1(n1123), .A2(n1082), .Y(n420) );
  NAND2X0_LVT U293 ( .A1(n1136), .A2(n1080), .Y(n497) );
  NAND4X0_LVT U294 ( .A1(n104), .A2(n119), .A3(n420), .A4(n497), .Y(n306) );
  AO22X1_LVT U295 ( .A1(n1087), .A2(n105), .A3(n985), .A4(n306), .Y(n106) );
  INVX1_LVT U296 ( .A(n106), .Y(n113) );
  AND2X1_LVT U297 ( .A1(n107), .A2(n1088), .Y(n109) );
  OR2X1_LVT U298 ( .A1(opv2[7]), .A2(n1126), .Y(n108) );
  NAND2X0_LVT U301 ( .A1(opv2[4]), .A2(n350), .Y(n805) );
  INVX1_LVT U302 ( .A(n805), .Y(n703) );
  NAND2X0_LVT U303 ( .A1(n1085), .A2(n1112), .Y(n411) );
  NAND2X0_LVT U304 ( .A1(n1121), .A2(n1082), .Y(n568) );
  NAND2X0_LVT U305 ( .A1(n1080), .A2(n1124), .Y(n1004) );
  NAND2X0_LVT U306 ( .A1(n1115), .A2(n16), .Y(n514) );
  NAND4X0_LVT U307 ( .A1(n411), .A2(n568), .A3(n1004), .A4(n514), .Y(n810) );
  MUX41X1_LVT U308 ( .A1(opv1[28]), .A3(opv1[27]), .A2(opv1[30]), .A4(opv1[29]), .S0(n1035), .S1(opv2[1]), .Y(n809) );
  AND2X1_LVT U309 ( .A1(n1085), .A2(n1143), .Y(n528) );
  AO222X1_LVT U310 ( .A1(n810), .A2(n28), .A3(n809), .A4(n1083), .A5(n528), 
        .A6(n15), .Y(n427) );
  NAND2X0_LVT U311 ( .A1(n703), .A2(n427), .Y(n111) );
  FADDX1_LVT U314 ( .A(opv1[7]), .B(n116), .CI(n115), .CO(n710), .S(n117) );
  NAND2X0_LVT U315 ( .A1(n52), .A2(n117), .Y(n123) );
  INVX1_LVT U316 ( .A(n776), .Y(n122) );
  MUX41X1_LVT U317 ( .A1(opv1[0]), .A3(opv1[1]), .A2(n1122), .A4(n1142), .S0(
        n1035), .S1(n1036), .Y(n867) );
  NAND2X0_LVT U318 ( .A1(n1125), .A2(n16), .Y(n255) );
  NAND2X0_LVT U319 ( .A1(n1080), .A2(n1114), .Y(n259) );
  NAND2X0_LVT U320 ( .A1(n1137), .A2(n1082), .Y(n307) );
  NAND4X0_LVT U321 ( .A1(n255), .A2(n259), .A3(n119), .A4(n307), .Y(n860) );
  AO22X1_LVT U322 ( .A1(n1083), .A2(n867), .A3(n28), .A4(n860), .Y(n438) );
  NAND2X0_LVT U323 ( .A1(n438), .A2(n1086), .Y(n121) );
  NAND2X0_LVT U324 ( .A1(n66), .A2(link_addr[7]), .Y(n120) );
  NAND2X0_LVT U327 ( .A1(n1133), .A2(n1082), .Y(n423) );
  NAND2X0_LVT U328 ( .A1(n1085), .A2(n1120), .Y(n416) );
  NAND2X0_LVT U329 ( .A1(n1127), .A2(n16), .Y(n493) );
  NAND2X0_LVT U330 ( .A1(n1130), .A2(n1080), .Y(n500) );
  NAND4X0_LVT U331 ( .A1(n423), .A2(n416), .A3(n493), .A4(n500), .Y(n804) );
  NAND2X0_LVT U332 ( .A1(n1085), .A2(n1135), .Y(n424) );
  NAND2X0_LVT U333 ( .A1(n1119), .A2(n1082), .Y(n410) );
  NAND2X0_LVT U334 ( .A1(n1128), .A2(n16), .Y(n501) );
  NAND2X0_LVT U335 ( .A1(n1113), .A2(n1080), .Y(n513) );
  NAND4X0_LVT U336 ( .A1(n424), .A2(n410), .A3(n501), .A4(n513), .Y(n811) );
  NAND2X0_LVT U337 ( .A1(n1085), .A2(n1132), .Y(n419) );
  NAND2X0_LVT U338 ( .A1(n1134), .A2(n1082), .Y(n415) );
  NAND2X0_LVT U339 ( .A1(n1116), .A2(n16), .Y(n496) );
  NAND2X0_LVT U340 ( .A1(n1117), .A2(n1080), .Y(n492) );
  NAND4X0_LVT U341 ( .A1(n419), .A2(n415), .A3(n496), .A4(n492), .Y(n731) );
  AO222X1_LVT U342 ( .A1(n804), .A2(n15), .A3(n811), .A4(n19), .A5(n731), .A6(
        n1083), .Y(n125) );
  NAND2X0_LVT U343 ( .A1(n1090), .A2(n125), .Y(n126) );
  NAND2X0_LVT U345 ( .A1(opv1[0]), .A2(mem_offset[0]), .Y(n605) );
  AND2X1_LVT U350 ( .A1(n605), .A2(n130), .Y(n132) );
  OR2X1_LVT U351 ( .A1(mem_offset[0]), .A2(opv1[0]), .Y(n131) );
  AND2X1_LVT U352 ( .A1(n132), .A2(n131), .Y(mem_addr[0]) );
  FADDX1_LVT U353 ( .A(n2), .B(opv1[0]), .CI(n133), .CO(n253), .S(n134) );
  NAND2X0_LVT U354 ( .A1(n52), .A2(n134), .Y(n252) );
  AO22X1_LVT U355 ( .A1(N287), .A2(n546), .A3(n1001), .A4(n1086), .Y(n241) );
  NAND2X0_LVT U356 ( .A1(n1085), .A2(n1128), .Y(n478) );
  NAND2X0_LVT U357 ( .A1(n1113), .A2(n1082), .Y(n450) );
  NAND4X0_LVT U358 ( .A1(n136), .A2(n135), .A3(n478), .A4(n450), .Y(n756) );
  NAND2X0_LVT U359 ( .A1(n1085), .A2(n1127), .Y(n470) );
  NAND2X0_LVT U360 ( .A1(n1130), .A2(n1082), .Y(n477) );
  NAND4X0_LVT U361 ( .A1(n138), .A2(n137), .A3(n470), .A4(n477), .Y(n758) );
  AO22X1_LVT U362 ( .A1(opv2[1]), .A2(n139), .A3(n1085), .A4(opv1[28]), .Y(
        n140) );
  AO21X1_LVT U363 ( .A1(opv1[29]), .A2(n16), .A3(n140), .Y(n742) );
  NAND2X0_LVT U364 ( .A1(opv1[26]), .A2(n1082), .Y(n539) );
  NAND2X0_LVT U365 ( .A1(n1085), .A2(n1115), .Y(n451) );
  NAND4X0_LVT U366 ( .A1(n142), .A2(n141), .A3(n539), .A4(n451), .Y(n757) );
  AO22X1_LVT U367 ( .A1(opv2[2]), .A2(n742), .A3(n1038), .A4(n757), .Y(n709)
         );
  AO222X1_LVT U368 ( .A1(n756), .A2(n1083), .A3(n758), .A4(n28), .A5(n709), 
        .A6(opv2[3]), .Y(n834) );
  NAND2X0_LVT U369 ( .A1(n1117), .A2(n1082), .Y(n469) );
  NAND2X0_LVT U370 ( .A1(n1085), .A2(n1116), .Y(n474) );
  NAND4X0_LVT U371 ( .A1(n144), .A2(n143), .A3(n469), .A4(n474), .Y(n743) );
  NAND2X0_LVT U372 ( .A1(n1085), .A2(n1129), .Y(n462) );
  NAND2X0_LVT U373 ( .A1(n1136), .A2(n1082), .Y(n473) );
  NAND4X0_LVT U374 ( .A1(n146), .A2(n145), .A3(n462), .A4(n473), .Y(n686) );
  AO22X1_LVT U375 ( .A1(opv2[2]), .A2(n743), .A3(n1038), .A4(n686), .Y(n718)
         );
  NAND2X0_LVT U376 ( .A1(n1085), .A2(n1114), .Y(n459) );
  NAND2X0_LVT U377 ( .A1(n1125), .A2(n1082), .Y(n463) );
  NAND4X0_LVT U378 ( .A1(n148), .A2(n147), .A3(n459), .A4(n463), .Y(n672) );
  AO22X1_LVT U379 ( .A1(opv2[3]), .A2(n718), .A3(n1084), .A4(n672), .Y(n154)
         );
  INVX1_LVT U380 ( .A(n587), .Y(n312) );
  NAND2X0_LVT U381 ( .A1(n1122), .A2(n1082), .Y(n458) );
  NAND3X0_LVT U382 ( .A1(n151), .A2(n150), .A3(n458), .Y(n152) );
  AO22X1_LVT U383 ( .A1(opv1[0]), .A2(n312), .A3(n311), .A4(n152), .Y(n153) );
  AO221X1_LVT U384 ( .A1(opv2[4]), .A2(n834), .A3(n1042), .A4(n154), .A5(n153), 
        .Y(n239) );
  NAND2X0_LVT U386 ( .A1(n1143), .A2(n1079), .Y(n155) );
  AND2X1_LVT U387 ( .A1(n155), .A2(n248), .Y(n237) );
  OA21X1_LVT U391 ( .A1(opv2[27]), .A2(n1070), .A3(opv2[26]), .Y(n156) );
  AO22X1_LVT U392 ( .A1(opv2[27]), .A2(n1070), .A3(n1071), .A4(n156), .Y(n227)
         );
  AO22X1_LVT U395 ( .A1(opv2[25]), .A2(n1073), .A3(opv2[24]), .A4(n1072), .Y(
        n225) );
  OR2X1_LVT U396 ( .A1(n1072), .A2(opv2[24]), .Y(n445) );
  OA22X1_LVT U400 ( .A1(opv2[17]), .A2(n1059), .A3(opv2[18]), .A4(n1061), .Y(
        n157) );
  OA21X1_LVT U401 ( .A1(opv2[19]), .A2(n1062), .A3(n157), .Y(n207) );
  AO22X1_LVT U403 ( .A1(opv2[16]), .A2(n1058), .A3(opv2[17]), .A4(n1059), .Y(
        n162) );
  NAND2X0_LVT U405 ( .A1(n1135), .A2(n1060), .Y(n161) );
  AO22X1_LVT U406 ( .A1(opv2[18]), .A2(n1061), .A3(opv2[19]), .A4(n1062), .Y(
        n160) );
  AO22X1_LVT U407 ( .A1(n207), .A2(n162), .A3(n161), .A4(n160), .Y(n208) );
  OA22X1_LVT U411 ( .A1(opv2[13]), .A2(n1054), .A3(opv2[14]), .A4(n1056), .Y(
        n163) );
  OA21X1_LVT U412 ( .A1(opv2[15]), .A2(n1057), .A3(n163), .Y(n194) );
  AO22X1_LVT U414 ( .A1(opv2[13]), .A2(n1054), .A3(opv2[12]), .A4(n1053), .Y(
        n168) );
  NAND2X0_LVT U416 ( .A1(n1120), .A2(n1055), .Y(n167) );
  AO22X1_LVT U417 ( .A1(opv2[14]), .A2(n1056), .A3(opv2[15]), .A4(n1057), .Y(
        n166) );
  AO22X1_LVT U418 ( .A1(n194), .A2(n168), .A3(n167), .A4(n166), .Y(n200) );
  OA22X1_LVT U422 ( .A1(opv2[9]), .A2(n1049), .A3(opv2[10]), .A4(n1051), .Y(
        n169) );
  OA21X1_LVT U423 ( .A1(opv2[11]), .A2(n1052), .A3(n169), .Y(n197) );
  AO22X1_LVT U425 ( .A1(opv2[8]), .A2(n1048), .A3(opv2[9]), .A4(n1049), .Y(
        n174) );
  NAND2X0_LVT U427 ( .A1(n1132), .A2(n1050), .Y(n173) );
  AO22X1_LVT U428 ( .A1(opv2[10]), .A2(n1051), .A3(opv2[11]), .A4(n1052), .Y(
        n172) );
  AO22X1_LVT U429 ( .A1(n197), .A2(n174), .A3(n173), .A4(n172), .Y(n198) );
  AO222X1_LVT U433 ( .A1(n1037), .A2(n1039), .A3(n1037), .A4(n1080), .A5(n1039), .A6(opv2[1]), .Y(n175) );
  AND2X1_LVT U434 ( .A1(n176), .A2(n175), .Y(n178) );
  OR2X1_LVT U435 ( .A1(n1041), .A2(opv2[2]), .Y(n177) );
  AND2X1_LVT U436 ( .A1(n178), .A2(n177), .Y(n181) );
  NAND2X0_LVT U437 ( .A1(n1142), .A2(n1040), .Y(n179) );
  OA221X1_LVT U438 ( .A1(n181), .A2(opv2[2]), .A3(n181), .A4(n1041), .A5(n179), 
        .Y(n182) );
  AO21X1_LVT U439 ( .A1(opv2[3]), .A2(n1043), .A3(n182), .Y(n184) );
  AO222X1_LVT U441 ( .A1(opv2[4]), .A2(n184), .A3(opv2[4]), .A4(n1044), .A5(
        n184), .A6(n1044), .Y(n185) );
  AO222X1_LVT U442 ( .A1(opv2[5]), .A2(n1045), .A3(opv2[5]), .A4(n185), .A5(
        n1045), .A6(n185), .Y(n188) );
  AO222X1_LVT U444 ( .A1(opv2[6]), .A2(n188), .A3(opv2[6]), .A4(n1046), .A5(
        n188), .A6(n1046), .Y(n192) );
  OA22X1_LVT U446 ( .A1(opv2[7]), .A2(n1047), .A3(opv2[8]), .A4(n1048), .Y(
        n190) );
  OA221X1_LVT U447 ( .A1(n192), .A2(opv2[7]), .A3(n192), .A4(n1047), .A5(n190), 
        .Y(n196) );
  AO22X1_LVT U448 ( .A1(n194), .A2(opv2[12]), .A3(n194), .A4(n1053), .Y(n195)
         );
  OA221X1_LVT U449 ( .A1(n198), .A2(n197), .A3(n198), .A4(n196), .A5(n195), 
        .Y(n199) );
  OA22X1_LVT U450 ( .A1(opv2[16]), .A2(n1058), .A3(n200), .A4(n199), .Y(n206)
         );
  OR2X1_LVT U452 ( .A1(n1065), .A2(opv2[21]), .Y(n202) );
  OA22X1_LVT U455 ( .A1(opv2[22]), .A2(n1067), .A3(opv2[23]), .A4(n1066), .Y(
        n216) );
  AND2X1_LVT U456 ( .A1(n202), .A2(n216), .Y(n204) );
  OR2X1_LVT U458 ( .A1(n1063), .A2(opv2[20]), .Y(n203) );
  AND2X1_LVT U459 ( .A1(n204), .A2(n203), .Y(n205) );
  OA221X1_LVT U460 ( .A1(n208), .A2(n207), .A3(n208), .A4(n206), .A5(n205), 
        .Y(n209) );
  INVX1_LVT U461 ( .A(n209), .Y(n219) );
  AND2X1_LVT U462 ( .A1(opv2[22]), .A2(n1067), .Y(n385) );
  OR2X1_LVT U463 ( .A1(n1066), .A2(opv2[23]), .Y(n408) );
  AO22X1_LVT U464 ( .A1(n385), .A2(n408), .A3(opv2[23]), .A4(n1066), .Y(n211)
         );
  INVX1_LVT U465 ( .A(n211), .Y(n218) );
  OA21X1_LVT U466 ( .A1(opv2[21]), .A2(n1065), .A3(opv2[20]), .Y(n212) );
  AO22X1_LVT U467 ( .A1(opv2[21]), .A2(n1065), .A3(n1063), .A4(n212), .Y(n215)
         );
  NAND2X0_LVT U468 ( .A1(n216), .A2(n215), .Y(n217) );
  NAND3X0_LVT U469 ( .A1(n219), .A2(n218), .A3(n217), .Y(n224) );
  NAND2X0_LVT U471 ( .A1(opv1[26]), .A2(n1069), .Y(n939) );
  NAND2X0_LVT U473 ( .A1(opv1[27]), .A2(n1068), .Y(n964) );
  AND2X1_LVT U474 ( .A1(n939), .A2(n964), .Y(n222) );
  OR2X1_LVT U475 ( .A1(n1073), .A2(opv2[25]), .Y(n221) );
  AND2X1_LVT U476 ( .A1(n222), .A2(n221), .Y(n223) );
  OA221X1_LVT U477 ( .A1(n225), .A2(n445), .A3(n225), .A4(n224), .A5(n223), 
        .Y(n226) );
  OAI22X1_LVT U479 ( .A1(n227), .A2(n226), .A3(opv2[28]), .A4(n1075), .Y(n229)
         );
  NAND2X0_LVT U480 ( .A1(opv2[28]), .A2(n1075), .Y(n552) );
  AO22X1_LVT U481 ( .A1(opv1[29]), .A2(n1077), .A3(n229), .A4(n552), .Y(n232)
         );
  AO221X1_LVT U482 ( .A1(n232), .A2(opv1[29]), .A3(n232), .A4(n1077), .A5(n230), .Y(n233) );
  NAND2X0_LVT U483 ( .A1(n234), .A2(n233), .Y(n245) );
  AND2X1_LVT U485 ( .A1(opv2[31]), .A2(n1074), .Y(n235) );
  OR2X1_LVT U486 ( .A1(n245), .A2(n235), .Y(n236) );
  AND2X1_LVT U487 ( .A1(n237), .A2(n236), .Y(n238) );
  AO22X1_LVT U488 ( .A1(n430), .A2(n239), .A3(n238), .A4(n1033), .Y(n240) );
  AOI22X1_LVT U489 ( .A1(opv1[0]), .A2(n241), .A3(aluop[1]), .A4(n240), .Y(
        n251) );
  AO222X1_LVT U490 ( .A1(N287), .A2(n1033), .A3(N287), .A4(n1037), .A5(opv1[0]), .A6(n1035), .Y(n244) );
  AOI22X1_LVT U491 ( .A1(n66), .A2(link_addr[0]), .A3(n1088), .A4(n244), .Y(
        n250) );
  AO222X1_LVT U492 ( .A1(n1143), .A2(n1079), .A3(n1143), .A4(n245), .A5(n1079), 
        .A6(n245), .Y(n247) );
  NAND4X0_LVT U493 ( .A1(ex_aluop[0]), .A2(n248), .A3(n247), .A4(n1034), .Y(
        n249) );
  FADDX1_LVT U495 ( .A(opv1[1]), .B(n254), .CI(n253), .CO(n279), .S(n278) );
  AO222X1_LVT U496 ( .A1(n785), .A2(n1084), .A3(n783), .A4(n28), .A5(n520), 
        .A6(opv2[3]), .Y(n849) );
  NAND2X0_LVT U497 ( .A1(n1085), .A2(n1137), .Y(n256) );
  NAND2X0_LVT U498 ( .A1(n1080), .A2(n1129), .Y(n421) );
  NAND4X0_LVT U499 ( .A1(n257), .A2(n256), .A3(n255), .A4(n421), .Y(n691) );
  AO222X1_LVT U500 ( .A1(n701), .A2(n15), .A3(n765), .A4(n19), .A5(n691), .A6(
        n1083), .Y(n264) );
  NAND2X0_LVT U501 ( .A1(n1142), .A2(n1082), .Y(n261) );
  NAND2X0_LVT U502 ( .A1(n1122), .A2(n16), .Y(n260) );
  NAND3X0_LVT U503 ( .A1(n261), .A2(n260), .A3(n259), .Y(n262) );
  AO22X1_LVT U504 ( .A1(opv1[1]), .A2(n312), .A3(n311), .A4(n262), .Y(n263) );
  AO221X1_LVT U505 ( .A1(opv2[4]), .A2(n849), .A3(n1042), .A4(n264), .A5(n263), 
        .Y(n276) );
  NAND3X0_LVT U506 ( .A1(n1031), .A2(opv2[1]), .A3(opv1[1]), .Y(n266) );
  INVX1_LVT U507 ( .A(n266), .Y(n274) );
  AND2X2_LVT U508 ( .A1(n1086), .A2(n28), .Y(n957) );
  AO22X1_LVT U509 ( .A1(n66), .A2(link_addr[1]), .A3(n957), .A4(n846), .Y(n265) );
  INVX1_LVT U510 ( .A(n265), .Y(n272) );
  AND2X1_LVT U511 ( .A1(n266), .A2(n1088), .Y(n268) );
  OR2X1_LVT U512 ( .A1(opv1[1]), .A2(opv2[1]), .Y(n267) );
  AND3X1_LVT U515 ( .A1(n950), .A2(n777), .A3(n904), .Y(n319) );
  NAND2X0_LVT U516 ( .A1(n319), .A2(n847), .Y(n270) );
  NAND3X0_LVT U517 ( .A1(n272), .A2(n1093), .A3(n270), .Y(n273) );
  AO21X1_LVT U518 ( .A1(n274), .A2(n1087), .A3(n273), .Y(n275) );
  AO21X1_LVT U519 ( .A1(n350), .A2(n276), .A3(n275), .Y(n277) );
  FADDX1_LVT U521 ( .A(opv1[2]), .B(n280), .CI(n279), .CO(n304), .S(n281) );
  NAND2X0_LVT U522 ( .A1(n52), .A2(n281), .Y(n303) );
  NAND3X0_LVT U523 ( .A1(n1031), .A2(opv2[2]), .A3(n1122), .Y(n284) );
  INVX1_LVT U524 ( .A(n284), .Y(n282) );
  NAND2X0_LVT U525 ( .A1(n282), .A2(n1087), .Y(n302) );
  INVX1_LVT U526 ( .A(n319), .Y(n301) );
  AND2X1_LVT U529 ( .A1(n284), .A2(n1088), .Y(n286) );
  OR2X1_LVT U530 ( .A1(n1122), .A2(opv2[2]), .Y(n285) );
  AO222X1_LVT U533 ( .A1(n349), .A2(n1083), .A3(n347), .A4(n28), .A5(n933), 
        .A6(opv2[3]), .Y(n375) );
  NAND2X0_LVT U534 ( .A1(n1126), .A2(n16), .Y(n461) );
  NAND2X0_LVT U535 ( .A1(n1123), .A2(n1080), .Y(n472) );
  NAND4X0_LVT U536 ( .A1(n289), .A2(n288), .A3(n461), .A4(n472), .Y(n327) );
  AO222X1_LVT U537 ( .A1(n334), .A2(n15), .A3(n346), .A4(n19), .A5(n327), .A6(
        n1083), .Y(n294) );
  NAND2X0_LVT U538 ( .A1(n1142), .A2(n16), .Y(n457) );
  NAND2X0_LVT U539 ( .A1(n1080), .A2(n1137), .Y(n460) );
  NAND3X0_LVT U540 ( .A1(n291), .A2(n457), .A3(n460), .Y(n292) );
  AO22X1_LVT U541 ( .A1(n1122), .A2(n312), .A3(n311), .A4(n292), .Y(n293) );
  AO221X1_LVT U542 ( .A1(opv2[4]), .A2(n375), .A3(n1042), .A4(n294), .A5(n293), 
        .Y(n295) );
  NAND2X0_LVT U543 ( .A1(n350), .A2(n295), .Y(n296) );
  FADDX1_LVT U547 ( .A(opv1[3]), .B(n305), .CI(n304), .CO(n674), .S(n324) );
  AO22X1_LVT U548 ( .A1(opv2[2]), .A2(n528), .A3(n1038), .A4(n809), .Y(n955)
         );
  AO222X1_LVT U549 ( .A1(n810), .A2(n1083), .A3(n811), .A4(n28), .A5(n955), 
        .A6(opv2[3]), .Y(n862) );
  AO222X1_LVT U550 ( .A1(n731), .A2(n15), .A3(n804), .A4(n19), .A5(n306), .A6(
        n1083), .Y(n314) );
  NAND2X0_LVT U551 ( .A1(n1114), .A2(n16), .Y(n308) );
  NAND3X0_LVT U552 ( .A1(n309), .A2(n308), .A3(n307), .Y(n310) );
  AO22X1_LVT U553 ( .A1(n1142), .A2(n312), .A3(n311), .A4(n310), .Y(n313) );
  AO221X1_LVT U554 ( .A1(opv2[4]), .A2(n862), .A3(n1042), .A4(n314), .A5(n313), 
        .Y(n322) );
  AO22X1_LVT U555 ( .A1(n66), .A2(link_addr[3]), .A3(n957), .A4(n867), .Y(n320) );
  OA21X1_LVT U557 ( .A1(opv2[3]), .A2(n1142), .A3(n1088), .Y(n317) );
  NAND3X0_LVT U558 ( .A1(n1031), .A2(opv2[3]), .A3(n1142), .Y(n316) );
  MUX21X1_LVT U559 ( .A1(n1087), .A2(n317), .S0(n316), .Y(n318) );
  OR3X1_LVT U560 ( .A1(n320), .A2(n319), .A3(n318), .Y(n321) );
  AO21X1_LVT U561 ( .A1(n322), .A2(n350), .A3(n321), .Y(n323) );
  FADDX1_LVT U563 ( .A(opv1[6]), .B(n326), .CI(n325), .CO(n115), .S(n343) );
  AO22X1_LVT U564 ( .A1(n66), .A2(link_addr[6]), .A3(n985), .A4(n327), .Y(n341) );
  AO222X1_LVT U565 ( .A1(n349), .A2(n28), .A3(n348), .A4(n1083), .A5(n351), 
        .A6(n15), .Y(n392) );
  NAND3X0_LVT U566 ( .A1(n1031), .A2(n1125), .A3(opv2[6]), .Y(n330) );
  INVX1_LVT U567 ( .A(n330), .Y(n328) );
  AND2X1_LVT U568 ( .A1(n1086), .A2(n1040), .Y(n673) );
  AO22X1_LVT U569 ( .A1(n1087), .A2(n328), .A3(n386), .A4(n673), .Y(n329) );
  INVX1_LVT U570 ( .A(n329), .Y(n338) );
  AND2X1_LVT U571 ( .A1(n330), .A2(n1088), .Y(n332) );
  OR2X1_LVT U572 ( .A1(opv2[6]), .A2(n1125), .Y(n331) );
  AO222X1_LVT U575 ( .A1(n346), .A2(n15), .A3(n347), .A4(n19), .A5(n334), .A6(
        n1083), .Y(n335) );
  NAND2X0_LVT U576 ( .A1(n1090), .A2(n335), .Y(n336) );
  NAND3X0_LVT U577 ( .A1(n338), .A2(n1091), .A3(n336), .Y(n339) );
  AO21X1_LVT U578 ( .A1(n392), .A2(n703), .A3(n339), .Y(n340) );
  OR3X1_LVT U579 ( .A1(n776), .A2(n341), .A3(n340), .Y(n342) );
  FADDX1_LVT U581 ( .A(opv1[14]), .B(n345), .CI(n344), .CO(n790), .S(n367) );
  AO22X1_LVT U582 ( .A1(n66), .A2(link_addr[14]), .A3(n985), .A4(n346), .Y(
        n365) );
  NAND2X0_LVT U583 ( .A1(n1143), .A2(n777), .Y(n851) );
  INVX1_LVT U584 ( .A(n851), .Y(n919) );
  AO222X1_LVT U585 ( .A1(n349), .A2(n15), .A3(n348), .A4(n19), .A5(n347), .A6(
        n1083), .Y(n363) );
  NAND3X0_LVT U586 ( .A1(n1031), .A2(n1117), .A3(opv2[14]), .Y(n354) );
  INVX1_LVT U587 ( .A(n354), .Y(n352) );
  AND3X1_LVT U588 ( .A1(opv2[4]), .A2(n28), .A3(n350), .Y(n764) );
  AO22X1_LVT U589 ( .A1(n1087), .A2(n352), .A3(n351), .A4(n764), .Y(n353) );
  INVX1_LVT U590 ( .A(n353), .Y(n361) );
  AND2X1_LVT U591 ( .A1(n354), .A2(n1088), .Y(n356) );
  OR2X1_LVT U592 ( .A1(opv2[14]), .A2(n1117), .Y(n355) );
  NAND2X0_LVT U595 ( .A1(n1086), .A2(n358), .Y(n359) );
  NAND3X0_LVT U596 ( .A1(n361), .A2(n1096), .A3(n359), .Y(n362) );
  AO21X1_LVT U597 ( .A1(n1090), .A2(n363), .A3(n362), .Y(n364) );
  OR3X1_LVT U598 ( .A1(n365), .A2(n919), .A3(n364), .Y(n366) );
  FADDX1_LVT U600 ( .A(opv1[18]), .B(n369), .CI(n368), .CO(n864), .S(n370) );
  NAND2X0_LVT U601 ( .A1(n52), .A2(n370), .Y(n382) );
  NAND3X0_LVT U602 ( .A1(ex_aluop[0]), .A2(n1130), .A3(opv2[18]), .Y(n371) );
  OA21X1_LVT U603 ( .A1(n1130), .A2(opv2[18]), .A3(n371), .Y(n372) );
  AO22X1_LVT U604 ( .A1(n66), .A2(link_addr[18]), .A3(n1088), .A4(n372), .Y(
        n379) );
  AND2X1_LVT U605 ( .A1(n28), .A2(n1013), .Y(n868) );
  AO22X1_LVT U606 ( .A1(n957), .A2(n946), .A3(n868), .A4(n373), .Y(n378) );
  AO222X1_LVT U607 ( .A1(n387), .A2(n15), .A3(n374), .A4(n19), .A5(n945), .A6(
        n1084), .Y(n376) );
  AO22X1_LVT U608 ( .A1(n1086), .A2(n376), .A3(n1090), .A4(n375), .Y(n377) );
  NOR4X1_LVT U609 ( .A1(n919), .A2(n379), .A3(n378), .A4(n377), .Y(n381) );
  NAND3X0_LVT U610 ( .A1(n950), .A2(n987), .A3(n904), .Y(n879) );
  NAND4X0_LVT U611 ( .A1(ex_aluop[0]), .A2(n1130), .A3(opv2[18]), .A4(n1087), 
        .Y(n380) );
  FADDX1_LVT U613 ( .A(n1113), .B(n384), .CI(n383), .CO(n406), .S(n405) );
  AO22X1_LVT U614 ( .A1(opv2[22]), .A2(n529), .A3(n385), .A4(n1088), .Y(n403)
         );
  NAND2X0_LVT U615 ( .A1(n386), .A2(n1040), .Y(n391) );
  MUX41X1_LVT U616 ( .A1(n387), .A3(n946), .A2(n945), .A4(n947), .S0(n1040), 
        .S1(n1038), .Y(n388) );
  INVX1_LVT U617 ( .A(n388), .Y(n390) );
  AO221X1_LVT U618 ( .A1(opv2[4]), .A2(n391), .A3(n1042), .A4(n390), .A5(n389), 
        .Y(n397) );
  NAND3X0_LVT U619 ( .A1(aluop[1]), .A2(n1042), .A3(n392), .Y(n396) );
  NAND2X0_LVT U620 ( .A1(n393), .A2(n1042), .Y(n394) );
  NAND3X0_LVT U621 ( .A1(n1139), .A2(n1143), .A3(n394), .Y(n395) );
  NAND3X0_LVT U622 ( .A1(n397), .A2(n396), .A3(n395), .Y(n400) );
  AO22X1_LVT U624 ( .A1(opv2[22]), .A2(n546), .A3(n1064), .A4(n1088), .Y(n399)
         );
  AO22X1_LVT U625 ( .A1(n430), .A2(n400), .A3(n1113), .A4(n399), .Y(n402) );
  AND2X1_LVT U626 ( .A1(n66), .A2(link_addr[22]), .Y(n401) );
  OR3X1_LVT U627 ( .A1(n403), .A2(n402), .A3(n401), .Y(n404) );
  FADDX1_LVT U629 ( .A(n1112), .B(n407), .CI(n406), .CO(n443), .S(n442) );
  INVX1_LVT U630 ( .A(n408), .Y(n440) );
  AO221X1_LVT U631 ( .A1(n1112), .A2(n546), .A3(n1066), .A4(n1088), .A5(n529), 
        .Y(n414) );
  NAND4X0_LVT U632 ( .A1(n413), .A2(n412), .A3(n411), .A4(n410), .Y(n963) );
  AOI22X1_LVT U633 ( .A1(opv2[23]), .A2(n414), .A3(n957), .A4(n963), .Y(n436)
         );
  NAND4X0_LVT U634 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .Y(n961) );
  NAND4X0_LVT U635 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .Y(n861) );
  NAND4X0_LVT U636 ( .A1(n426), .A2(n425), .A3(n424), .A4(n423), .Y(n962) );
  AO222X1_LVT U637 ( .A1(n961), .A2(n15), .A3(n861), .A4(n19), .A5(n962), .A6(
        n1083), .Y(n428) );
  AOI22X1_LVT U638 ( .A1(n1086), .A2(n428), .A3(n1090), .A4(n427), .Y(n435) );
  NAND2X0_LVT U639 ( .A1(n430), .A2(n1139), .Y(n585) );
  INVX1_LVT U640 ( .A(n585), .Y(n433) );
  NAND2X0_LVT U642 ( .A1(n1040), .A2(n1042), .Y(n431) );
  NAND3X0_LVT U643 ( .A1(n433), .A2(n1143), .A3(n431), .Y(n970) );
  NAND2X0_LVT U644 ( .A1(n66), .A2(link_addr[23]), .Y(n434) );
  NAND4X0_LVT U645 ( .A1(n436), .A2(n435), .A3(n970), .A4(n434), .Y(n437) );
  AO21X1_LVT U646 ( .A1(n438), .A2(n1013), .A3(n437), .Y(n439) );
  AO21X1_LVT U647 ( .A1(n1088), .A2(n440), .A3(n439), .Y(n441) );
  FADDX1_LVT U649 ( .A(n1115), .B(n444), .CI(n443), .CO(n488), .S(n487) );
  AND2X1_LVT U650 ( .A1(n1090), .A2(n1040), .Y(n954) );
  AO22X1_LVT U651 ( .A1(n709), .A2(n954), .A3(n987), .A4(n708), .Y(n485) );
  INVX1_LVT U652 ( .A(n445), .Y(n446) );
  AO22X1_LVT U653 ( .A1(n446), .A2(n1088), .A3(n66), .A4(link_addr[24]), .Y(
        n447) );
  INVX1_LVT U654 ( .A(n447), .Y(n454) );
  INVX1_LVT U655 ( .A(n919), .Y(n453) );
  NAND4X0_LVT U656 ( .A1(n451), .A2(n450), .A3(n449), .A4(n448), .Y(n534) );
  NAND2X0_LVT U657 ( .A1(n957), .A2(n534), .Y(n452) );
  NAND3X0_LVT U658 ( .A1(n454), .A2(n453), .A3(n452), .Y(n484) );
  NAND2X0_LVT U659 ( .A1(opv1[1]), .A2(n1080), .Y(n456) );
  NAND4X0_LVT U660 ( .A1(n459), .A2(n458), .A3(n457), .A4(n456), .Y(n829) );
  NAND4X0_LVT U661 ( .A1(n463), .A2(n462), .A3(n461), .A4(n460), .Y(n891) );
  AO22X1_LVT U662 ( .A1(n1084), .A2(n829), .A3(n28), .A4(n891), .Y(n466) );
  INVX1_LVT U663 ( .A(n464), .Y(n465) );
  OA222X1_LVT U664 ( .A1(n466), .A2(opv1[0]), .A3(n466), .A4(opv2[3]), .A5(
        n466), .A6(n465), .Y(n720) );
  NAND4X0_LVT U665 ( .A1(n470), .A2(n469), .A3(n468), .A4(n467), .Y(n890) );
  NAND4X0_LVT U666 ( .A1(n474), .A2(n473), .A3(n472), .A4(n471), .Y(n892) );
  NAND4X0_LVT U667 ( .A1(n478), .A2(n477), .A3(n476), .A4(n475), .Y(n886) );
  AO222X1_LVT U668 ( .A1(n890), .A2(n15), .A3(n892), .A4(n19), .A5(n886), .A6(
        n1084), .Y(n481) );
  AO221X1_LVT U669 ( .A1(n1115), .A2(n546), .A3(n1072), .A4(n1088), .A5(n529), 
        .Y(n480) );
  AO22X1_LVT U670 ( .A1(n1086), .A2(n481), .A3(opv2[24]), .A4(n480), .Y(n482)
         );
  AO21X1_LVT U671 ( .A1(n720), .A2(n1013), .A3(n482), .Y(n483) );
  OR3X1_LVT U672 ( .A1(n485), .A2(n484), .A3(n483), .Y(n486) );
  FADDX1_LVT U674 ( .A(n1121), .B(n489), .CI(n488), .CO(n935), .S(n525) );
  NAND3X0_LVT U675 ( .A1(n1031), .A2(n1121), .A3(opv2[25]), .Y(n507) );
  AND2X1_LVT U676 ( .A1(n507), .A2(n1088), .Y(n491) );
  OR2X1_LVT U677 ( .A1(opv2[25]), .A2(n1121), .Y(n490) );
  AND2X1_LVT U678 ( .A1(n491), .A2(n490), .Y(n523) );
  NAND4X0_LVT U679 ( .A1(n495), .A2(n494), .A3(n493), .A4(n492), .Y(n999) );
  NAND4X0_LVT U680 ( .A1(n499), .A2(n498), .A3(n497), .A4(n496), .Y(n925) );
  NAND4X0_LVT U681 ( .A1(n503), .A2(n502), .A3(n501), .A4(n500), .Y(n994) );
  AO222X1_LVT U682 ( .A1(n999), .A2(n15), .A3(n925), .A4(n19), .A5(n994), .A6(
        n1083), .Y(n505) );
  INVX1_LVT U685 ( .A(n987), .Y(n508) );
  OA22X1_LVT U686 ( .A1(n509), .A2(n508), .A3(n798), .A4(n507), .Y(n511) );
  NAND2X0_LVT U687 ( .A1(link_addr[25]), .A2(n66), .Y(n510) );
  NAND4X0_LVT U690 ( .A1(n516), .A2(n515), .A3(n514), .A4(n513), .Y(n996) );
  NAND2X0_LVT U691 ( .A1(n957), .A2(n996), .Y(n517) );
  NAND3X0_LVT U692 ( .A1(n1098), .A2(n1097), .A3(n517), .Y(n522) );
  AND2X1_LVT U693 ( .A1(n954), .A2(n520), .Y(n521) );
  OR3X1_LVT U694 ( .A1(n523), .A2(n522), .A3(n521), .Y(n524) );
  FADDX1_LVT U696 ( .A(n1140), .B(n527), .CI(n526), .CO(n988), .S(n558) );
  OR2X1_LVT U697 ( .A1(n950), .A2(n528), .Y(n900) );
  AO22X1_LVT U698 ( .A1(opv2[28]), .A2(n529), .A3(n987), .A4(n900), .Y(n530)
         );
  INVX1_LVT U699 ( .A(n530), .Y(n533) );
  INVX1_LVT U700 ( .A(n970), .Y(n1019) );
  INVX1_LVT U701 ( .A(n1019), .Y(n532) );
  NAND2X0_LVT U702 ( .A1(n66), .A2(link_addr[28]), .Y(n531) );
  NAND3X0_LVT U703 ( .A1(n533), .A2(n532), .A3(n531), .Y(n556) );
  AO22X1_LVT U704 ( .A1(n1084), .A2(n534), .A3(n15), .A4(n886), .Y(n535) );
  INVX1_LVT U705 ( .A(n535), .Y(n543) );
  AO22X1_LVT U706 ( .A1(n1001), .A2(n1140), .A3(n19), .A4(n890), .Y(n536) );
  INVX1_LVT U707 ( .A(n536), .Y(n542) );
  NAND2X0_LVT U708 ( .A1(n1141), .A2(n16), .Y(n538) );
  NAND3X0_LVT U709 ( .A1(n539), .A2(n538), .A3(n537), .Y(n540) );
  NAND2X0_LVT U710 ( .A1(n28), .A2(n540), .Y(n541) );
  NAND3X0_LVT U711 ( .A1(n543), .A2(n542), .A3(n541), .Y(n544) );
  OA222X1_LVT U712 ( .A1(n1038), .A2(n1085), .A3(n1038), .A4(opv1[0]), .A5(
        opv2[2]), .A6(n829), .Y(n899) );
  AO222X1_LVT U713 ( .A1(n891), .A2(n1083), .A3(n892), .A4(n28), .A5(n899), 
        .A6(opv2[3]), .Y(n760) );
  AO22X1_LVT U714 ( .A1(n1086), .A2(n544), .A3(n1013), .A4(n760), .Y(n545) );
  INVX1_LVT U715 ( .A(n545), .Y(n551) );
  OA221X1_LVT U717 ( .A1(opv2[28]), .A2(n1088), .A3(n1076), .A4(n546), .A5(
        n1140), .Y(n548) );
  INVX1_LVT U718 ( .A(n548), .Y(n550) );
  NAND2X0_LVT U719 ( .A1(n985), .A2(n742), .Y(n549) );
  NAND3X0_LVT U720 ( .A1(n551), .A2(n550), .A3(n549), .Y(n555) );
  INVX1_LVT U721 ( .A(n552), .Y(n553) );
  AND2X1_LVT U722 ( .A1(n1088), .A2(n553), .Y(n554) );
  OR3X1_LVT U723 ( .A1(n556), .A2(n555), .A3(n554), .Y(n557) );
  FADDX1_LVT U725 ( .A(n1131), .B(n560), .CI(n559), .CO(n564), .S(n35) );
  XOR2X1_LVT U726 ( .A1(n1139), .A2(opv2[31]), .Y(n562) );
  XOR2X1_LVT U727 ( .A1(n562), .A2(n1143), .Y(n563) );
  XOR2X1_LVT U728 ( .A1(n564), .A2(n563), .Y(n602) );
  NAND2X0_LVT U729 ( .A1(n66), .A2(link_addr[31]), .Y(n600) );
  NAND3X0_LVT U730 ( .A1(ex_aluop[0]), .A2(n1143), .A3(opv2[31]), .Y(n565) );
  NAND2X0_LVT U731 ( .A1(n1088), .A2(n565), .Y(n586) );
  OA22X1_LVT U732 ( .A1(n1079), .A2(n586), .A3(n798), .A4(n565), .Y(n599) );
  NAND2X0_LVT U733 ( .A1(n1085), .A2(n1141), .Y(n569) );
  NAND4X0_LVT U734 ( .A1(n571), .A2(n570), .A3(n569), .A4(n568), .Y(n956) );
  NAND2X0_LVT U735 ( .A1(opv1[29]), .A2(n1082), .Y(n573) );
  NAND3X0_LVT U736 ( .A1(n575), .A2(n574), .A3(n573), .Y(n576) );
  AO22X1_LVT U737 ( .A1(n1084), .A2(n956), .A3(n28), .A4(n576), .Y(n577) );
  INVX1_LVT U738 ( .A(n577), .Y(n583) );
  AO22X1_LVT U740 ( .A1(n1001), .A2(n1143), .A3(n19), .A4(n962), .Y(n580) );
  INVX1_LVT U741 ( .A(n580), .Y(n582) );
  NAND2X0_LVT U742 ( .A1(n15), .A2(n963), .Y(n581) );
  NAND3X0_LVT U743 ( .A1(n583), .A2(n582), .A3(n581), .Y(n584) );
  NAND2X0_LVT U744 ( .A1(n1086), .A2(n584), .Y(n598) );
  AND2X1_LVT U745 ( .A1(n586), .A2(n585), .Y(n592) );
  INVX1_LVT U746 ( .A(n587), .Y(n590) );
  INVX1_LVT U747 ( .A(n588), .Y(n589) );
  NAND2X0_LVT U748 ( .A1(n590), .A2(n589), .Y(n591) );
  AND2X1_LVT U749 ( .A1(n592), .A2(n591), .Y(n596) );
  MUX41X1_LVT U750 ( .A1(n867), .A3(n861), .A2(n860), .A4(n961), .S0(n1040), 
        .S1(n1038), .Y(n594) );
  INVX1_LVT U751 ( .A(n594), .Y(n814) );
  OA22X1_LVT U752 ( .A1(n596), .A2(n1074), .A3(n814), .A4(n976), .Y(n597) );
  NAND4X0_LVT U753 ( .A1(n600), .A2(n599), .A3(n598), .A4(n597), .Y(n601) );
  FADDX1_LVT U756 ( .A(mem_offset[1]), .B(n1039), .CI(n605), .S(n604) );
  AND2X1_LVT U757 ( .A1(n130), .A2(n604), .Y(mem_addr[1]) );
  INVX1_LVT U758 ( .A(n605), .Y(n606) );
  AO222X1_LVT U759 ( .A1(opv1[1]), .A2(n606), .A3(opv1[1]), .A4(mem_offset[1]), 
        .A5(n606), .A6(mem_offset[1]), .Y(n608) );
  AND2X1_LVT U760 ( .A1(n130), .A2(n607), .Y(mem_addr[2]) );
  FADDX1_LVT U761 ( .A(opv1[2]), .B(mem_offset[2]), .CI(n608), .CO(n610), .S(
        n607) );
  AND2X1_LVT U762 ( .A1(n130), .A2(n609), .Y(mem_addr[3]) );
  FADDX1_LVT U763 ( .A(opv1[3]), .B(mem_offset[3]), .CI(n610), .CO(n612), .S(
        n609) );
  AND2X1_LVT U764 ( .A1(n130), .A2(n611), .Y(mem_addr[4]) );
  FADDX1_LVT U765 ( .A(n1114), .B(mem_offset[4]), .CI(n612), .CO(n614), .S(
        n611) );
  AND2X1_LVT U766 ( .A1(n130), .A2(n613), .Y(mem_addr[5]) );
  FADDX1_LVT U767 ( .A(opv1[5]), .B(mem_offset[5]), .CI(n614), .CO(n616), .S(
        n613) );
  AND2X1_LVT U768 ( .A1(n130), .A2(n615), .Y(mem_addr[6]) );
  FADDX1_LVT U769 ( .A(opv1[6]), .B(mem_offset[6]), .CI(n616), .CO(n618), .S(
        n615) );
  AND2X1_LVT U770 ( .A1(n130), .A2(n617), .Y(mem_addr[7]) );
  FADDX1_LVT U771 ( .A(opv1[7]), .B(mem_offset[7]), .CI(n618), .CO(n620), .S(
        n617) );
  AND2X1_LVT U772 ( .A1(n130), .A2(n619), .Y(mem_addr[8]) );
  FADDX1_LVT U773 ( .A(opv1[8]), .B(mem_offset[8]), .CI(n620), .CO(n622), .S(
        n619) );
  AND2X1_LVT U774 ( .A1(n130), .A2(n621), .Y(mem_addr[9]) );
  FADDX1_LVT U775 ( .A(opv1[9]), .B(mem_offset[9]), .CI(n622), .CO(n624), .S(
        n621) );
  AND2X1_LVT U776 ( .A1(n130), .A2(n623), .Y(mem_addr[10]) );
  FADDX1_LVT U777 ( .A(opv1[10]), .B(mem_offset[10]), .CI(n624), .CO(n626), 
        .S(n623) );
  AND2X1_LVT U778 ( .A1(n130), .A2(n625), .Y(mem_addr[11]) );
  FADDX1_LVT U779 ( .A(opv1[11]), .B(mem_offset[11]), .CI(n626), .CO(n628), 
        .S(n625) );
  AND2X1_LVT U780 ( .A1(n130), .A2(n627), .Y(mem_addr[12]) );
  FADDX1_LVT U781 ( .A(n1116), .B(mem_offset[12]), .CI(n628), .CO(n630), .S(
        n627) );
  AND2X1_LVT U782 ( .A1(n130), .A2(n629), .Y(mem_addr[13]) );
  FADDX1_LVT U783 ( .A(opv1[13]), .B(mem_offset[13]), .CI(n630), .CO(n633), 
        .S(n629) );
  AND2X1_LVT U784 ( .A1(n130), .A2(n631), .Y(mem_addr[14]) );
  FADDX1_LVT U786 ( .A(n1117), .B(mem_offset[14]), .CI(n633), .CO(n635), .S(
        n631) );
  AND2X1_LVT U787 ( .A1(n130), .A2(n634), .Y(mem_addr[15]) );
  FADDX1_LVT U788 ( .A(n1120), .B(mem_offset[15]), .CI(n635), .CO(n637), .S(
        n634) );
  AND2X1_LVT U789 ( .A1(n130), .A2(n636), .Y(mem_addr[16]) );
  FADDX1_LVT U790 ( .A(opv1[16]), .B(mem_offset[16]), .CI(n637), .CO(n639), 
        .S(n636) );
  AND2X1_LVT U791 ( .A1(n130), .A2(n638), .Y(mem_addr[17]) );
  FADDX1_LVT U792 ( .A(opv1[17]), .B(mem_offset[17]), .CI(n639), .CO(n641), 
        .S(n638) );
  AND2X1_LVT U793 ( .A1(n130), .A2(n640), .Y(mem_addr[18]) );
  FADDX1_LVT U794 ( .A(opv1[18]), .B(mem_offset[18]), .CI(n641), .CO(n643), 
        .S(n640) );
  AND2X1_LVT U795 ( .A1(n130), .A2(n642), .Y(mem_addr[19]) );
  FADDX1_LVT U796 ( .A(opv1[19]), .B(mem_offset[19]), .CI(n643), .CO(n645), 
        .S(n642) );
  AND2X1_LVT U797 ( .A1(n1144), .A2(n644), .Y(mem_addr[20]) );
  FADDX1_LVT U798 ( .A(opv1[20]), .B(mem_offset[20]), .CI(n645), .CO(n647), 
        .S(n644) );
  AND2X1_LVT U799 ( .A1(n130), .A2(n646), .Y(mem_addr[21]) );
  FADDX1_LVT U800 ( .A(n1119), .B(mem_offset[21]), .CI(n647), .CO(n649), .S(
        n646) );
  AND2X1_LVT U801 ( .A1(n1144), .A2(n648), .Y(mem_addr[22]) );
  FADDX1_LVT U802 ( .A(n1113), .B(mem_offset[22]), .CI(n649), .CO(n652), .S(
        n648) );
  AND2X1_LVT U803 ( .A1(n130), .A2(n650), .Y(mem_addr[23]) );
  FADDX1_LVT U804 ( .A(n1112), .B(mem_offset[23]), .CI(n652), .CO(n654), .S(
        n650) );
  AND2X1_LVT U805 ( .A1(n1144), .A2(n653), .Y(mem_addr[24]) );
  FADDX1_LVT U806 ( .A(n1115), .B(mem_offset[24]), .CI(n654), .CO(n656), .S(
        n653) );
  AND2X1_LVT U807 ( .A1(n130), .A2(n655), .Y(mem_addr[25]) );
  FADDX1_LVT U808 ( .A(n1121), .B(mem_offset[25]), .CI(n656), .CO(n658), .S(
        n655) );
  AND2X1_LVT U809 ( .A1(n130), .A2(n657), .Y(mem_addr[26]) );
  FADDX1_LVT U810 ( .A(n1124), .B(mem_offset[26]), .CI(n658), .CO(n660), .S(
        n657) );
  AND2X1_LVT U811 ( .A1(n130), .A2(n659), .Y(mem_addr[27]) );
  FADDX1_LVT U812 ( .A(n1141), .B(mem_offset[27]), .CI(n660), .CO(n662), .S(
        n659) );
  AND2X1_LVT U813 ( .A1(n1144), .A2(n661), .Y(mem_addr[28]) );
  FADDX1_LVT U814 ( .A(n1140), .B(mem_offset[28]), .CI(n662), .CO(n664), .S(
        n661) );
  AND2X1_LVT U815 ( .A1(n1144), .A2(n663), .Y(mem_addr[29]) );
  FADDX1_LVT U816 ( .A(opv1[29]), .B(mem_offset[29]), .CI(n664), .CO(n667), 
        .S(n663) );
  AND2X1_LVT U817 ( .A1(n1144), .A2(n665), .Y(mem_addr[30]) );
  FADDX1_LVT U818 ( .A(n1131), .B(mem_offset[30]), .CI(n667), .CO(n669), .S(
        n665) );
  XOR2X1_LVT U819 ( .A1(n1143), .A2(mem_offset[31]), .Y(n668) );
  XOR2X1_LVT U820 ( .A1(n669), .A2(n668), .Y(n671) );
  AND2X1_LVT U821 ( .A1(n671), .A2(n1144), .Y(mem_addr[31]) );
  AO22X1_LVT U822 ( .A1(n673), .A2(n899), .A3(n985), .A4(n672), .Y(n690) );
  FADDX1_LVT U823 ( .A(opv1[4]), .B(n675), .CI(n674), .CO(n692), .S(n685) );
  NAND2X0_LVT U824 ( .A1(n66), .A2(link_addr[4]), .Y(n683) );
  NAND4X0_LVT U825 ( .A1(n1031), .A2(opv2[4]), .A3(n1114), .A4(n1087), .Y(n682) );
  NAND3X0_LVT U826 ( .A1(n777), .A2(n904), .A3(n900), .Y(n681) );
  NAND2X0_LVT U827 ( .A1(n1044), .A2(n1042), .Y(n679) );
  NAND3X0_LVT U828 ( .A1(n1031), .A2(opv2[4]), .A3(n1114), .Y(n678) );
  NAND3X0_LVT U829 ( .A1(n1088), .A2(n679), .A3(n678), .Y(n680) );
  NAND4X0_LVT U830 ( .A1(n683), .A2(n682), .A3(n681), .A4(n680), .Y(n684) );
  AO21X1_LVT U831 ( .A1(n52), .A2(n685), .A3(n684), .Y(n689) );
  AO222X1_LVT U832 ( .A1(n758), .A2(n19), .A3(n743), .A4(n15), .A5(n686), .A6(
        n1084), .Y(n687) );
  AO222X1_LVT U833 ( .A1(n742), .A2(n15), .A3(n757), .A4(n1083), .A5(n756), 
        .A6(n28), .Y(n893) );
  AO22X1_LVT U834 ( .A1(n1090), .A2(n687), .A3(n703), .A4(n893), .Y(n688) );
  AO22X1_LVT U836 ( .A1(n1083), .A2(n846), .A3(n28), .A4(n839), .Y(n905) );
  AO22X1_LVT U837 ( .A1(n1086), .A2(n905), .A3(n985), .A4(n691), .Y(n707) );
  FADDX1_LVT U838 ( .A(opv1[5]), .B(n693), .CI(n692), .CO(n325), .S(n700) );
  AO21X1_LVT U839 ( .A1(n1143), .A2(n847), .A3(n950), .Y(n986) );
  AND2X1_LVT U840 ( .A1(n777), .A2(n904), .Y(n698) );
  OA21X1_LVT U841 ( .A1(n1137), .A2(opv2[5]), .A3(n1088), .Y(n695) );
  NAND3X0_LVT U842 ( .A1(n1031), .A2(n1137), .A3(opv2[5]), .Y(n694) );
  MUX21X1_LVT U843 ( .A1(n1087), .A2(n695), .S0(n694), .Y(n696) );
  AO21X1_LVT U844 ( .A1(n66), .A2(link_addr[5]), .A3(n696), .Y(n697) );
  AO21X1_LVT U845 ( .A1(n986), .A2(n698), .A3(n697), .Y(n699) );
  AO21X1_LVT U846 ( .A1(n52), .A2(n700), .A3(n699), .Y(n706) );
  AO222X1_LVT U847 ( .A1(n765), .A2(n15), .A3(n783), .A4(n19), .A5(n701), .A6(
        n1083), .Y(n704) );
  AO222X1_LVT U848 ( .A1(n785), .A2(n28), .A3(n984), .A4(n15), .A5(n784), .A6(
        n1083), .Y(n927) );
  AO22X1_LVT U849 ( .A1(n1090), .A2(n704), .A3(n703), .A4(n927), .Y(n705) );
  AO22X1_LVT U851 ( .A1(n709), .A2(n732), .A3(n777), .A4(n708), .Y(n723) );
  FADDX1_LVT U852 ( .A(opv1[8]), .B(n711), .CI(n710), .CO(n91), .S(n717) );
  OA21X1_LVT U853 ( .A1(n1129), .A2(opv2[8]), .A3(n1088), .Y(n715) );
  NAND3X0_LVT U854 ( .A1(n1031), .A2(n1129), .A3(opv2[8]), .Y(n714) );
  INVX1_LVT U855 ( .A(n714), .Y(n712) );
  AO22X1_LVT U856 ( .A1(n1087), .A2(n712), .A3(n66), .A4(link_addr[8]), .Y(
        n713) );
  AO21X1_LVT U857 ( .A1(n715), .A2(n714), .A3(n713), .Y(n716) );
  AO21X1_LVT U858 ( .A1(n52), .A2(n717), .A3(n716), .Y(n722) );
  AO222X1_LVT U859 ( .A1(n1040), .A2(n718), .A3(n756), .A4(n19), .A5(n758), 
        .A6(n15), .Y(n719) );
  AO22X1_LVT U860 ( .A1(n1086), .A2(n720), .A3(n1090), .A4(n719), .Y(n721) );
  AO222X1_LVT U862 ( .A1(n1132), .A2(n1033), .A3(n1132), .A4(n1050), .A5(
        opv2[11]), .A6(n1052), .Y(n727) );
  AO22X1_LVT U863 ( .A1(n66), .A2(link_addr[11]), .A3(n1088), .A4(n727), .Y(
        n738) );
  FADDX1_LVT U864 ( .A(opv1[11]), .B(n729), .CI(n728), .CO(n744), .S(n730) );
  AND2X1_LVT U865 ( .A1(n52), .A2(n730), .Y(n736) );
  AND3X1_LVT U866 ( .A1(ex_aluop[0]), .A2(n1132), .A3(opv2[11]), .Y(n734) );
  AO22X1_LVT U867 ( .A1(n955), .A2(n732), .A3(n985), .A4(n731), .Y(n733) );
  AO21X1_LVT U868 ( .A1(n734), .A2(n1087), .A3(n733), .Y(n735) );
  NOR4X1_LVT U869 ( .A1(n738), .A2(n737), .A3(n736), .A4(n735), .Y(n741) );
  AOI222X1_LVT U870 ( .A1(n860), .A2(n1083), .A3(n861), .A4(n28), .A5(n867), 
        .A6(n15), .Y(n977) );
  AOI222X1_LVT U871 ( .A1(n804), .A2(n1083), .A3(n811), .A4(n15), .A5(n810), 
        .A6(n19), .Y(n739) );
  OA22X1_LVT U872 ( .A1(n977), .A2(n1118), .A3(n739), .A4(n812), .Y(n740) );
  AO22X1_LVT U874 ( .A1(n985), .A2(n743), .A3(n764), .A4(n742), .Y(n763) );
  FADDX1_LVT U875 ( .A(opv1[12]), .B(n745), .CI(n744), .CO(n766), .S(n751) );
  OA21X1_LVT U876 ( .A1(n1116), .A2(opv2[12]), .A3(n1088), .Y(n749) );
  NAND3X0_LVT U877 ( .A1(ex_aluop[0]), .A2(n1116), .A3(opv2[12]), .Y(n748) );
  INVX1_LVT U878 ( .A(n748), .Y(n746) );
  AO22X1_LVT U879 ( .A1(n1087), .A2(n746), .A3(n66), .A4(link_addr[12]), .Y(
        n747) );
  AO21X1_LVT U880 ( .A1(n749), .A2(n748), .A3(n747), .Y(n750) );
  INVX1_LVT U883 ( .A(n776), .Y(n754) );
  NAND2X0_LVT U884 ( .A1(n777), .A2(n900), .Y(n753) );
  NAND3X0_LVT U885 ( .A1(n1105), .A2(n754), .A3(n753), .Y(n762) );
  AO222X1_LVT U886 ( .A1(n758), .A2(n1084), .A3(n757), .A4(n19), .A5(n756), 
        .A6(n15), .Y(n759) );
  AO22X1_LVT U887 ( .A1(n1086), .A2(n760), .A3(n1090), .A4(n759), .Y(n761) );
  AO22X1_LVT U889 ( .A1(n985), .A2(n765), .A3(n764), .A4(n984), .Y(n789) );
  FADDX1_LVT U890 ( .A(opv1[13]), .B(n767), .CI(n766), .CO(n344), .S(n774) );
  OA21X1_LVT U891 ( .A1(n1134), .A2(opv2[13]), .A3(n1088), .Y(n772) );
  NAND3X0_LVT U892 ( .A1(n1031), .A2(n1134), .A3(opv2[13]), .Y(n771) );
  INVX1_LVT U893 ( .A(n771), .Y(n769) );
  AO22X1_LVT U894 ( .A1(n1087), .A2(n769), .A3(n66), .A4(link_addr[13]), .Y(
        n770) );
  AO21X1_LVT U895 ( .A1(n772), .A2(n771), .A3(n770), .Y(n773) );
  INVX1_LVT U898 ( .A(n776), .Y(n779) );
  NAND2X0_LVT U899 ( .A1(n777), .A2(n986), .Y(n778) );
  NAND3X0_LVT U900 ( .A1(n1104), .A2(n779), .A3(n778), .Y(n788) );
  AO22X1_LVT U901 ( .A1(n1084), .A2(n926), .A3(n28), .A4(n925), .Y(n782) );
  AO22X1_LVT U902 ( .A1(n15), .A2(n839), .A3(n19), .A4(n846), .Y(n781) );
  OR2X1_LVT U903 ( .A1(n782), .A2(n781), .Y(n1012) );
  AO222X1_LVT U904 ( .A1(n785), .A2(n15), .A3(n784), .A4(n19), .A5(n783), .A6(
        n1083), .Y(n786) );
  AO22X1_LVT U905 ( .A1(n1086), .A2(n1012), .A3(n1090), .A4(n786), .Y(n787) );
  FADDX1_LVT U907 ( .A(opv1[15]), .B(n791), .CI(n790), .CO(n818), .S(n792) );
  NAND2X0_LVT U908 ( .A1(n52), .A2(n792), .Y(n803) );
  NAND3X0_LVT U909 ( .A1(ex_aluop[0]), .A2(n1120), .A3(opv2[15]), .Y(n799) );
  INVX1_LVT U910 ( .A(n799), .Y(n797) );
  AO21X1_LVT U911 ( .A1(n1057), .A2(n1055), .A3(n975), .Y(n796) );
  OR2X1_LVT U912 ( .A1(n797), .A2(n796), .Y(n802) );
  OR2X1_LVT U913 ( .A1(n799), .A2(n798), .Y(n801) );
  NAND2X0_LVT U914 ( .A1(n66), .A2(link_addr[15]), .Y(n800) );
  AND4X1_LVT U915 ( .A1(n803), .A2(n802), .A3(n801), .A4(n800), .Y(n817) );
  INVX1_LVT U916 ( .A(n804), .Y(n808) );
  NAND2X0_LVT U917 ( .A1(n1001), .A2(n1143), .Y(n806) );
  OA22X1_LVT U918 ( .A1(n808), .A2(n807), .A3(n806), .A4(n805), .Y(n816) );
  AOI222X1_LVT U919 ( .A1(n811), .A2(n1083), .A3(n810), .A4(n15), .A5(n809), 
        .A6(n19), .Y(n813) );
  OA22X1_LVT U920 ( .A1(n814), .A2(n1118), .A3(n813), .A4(n812), .Y(n815) );
  FADDX1_LVT U922 ( .A(opv1[16]), .B(n819), .CI(n818), .CO(n844), .S(n820) );
  NAND2X0_LVT U923 ( .A1(n52), .A2(n820), .Y(n823) );
  NAND4X0_LVT U924 ( .A1(n1031), .A2(n1127), .A3(opv2[16]), .A4(n1087), .Y(
        n822) );
  NAND3X0_LVT U925 ( .A1(opv1[0]), .A2(n1001), .A3(n1013), .Y(n821) );
  NAND4X0_LVT U926 ( .A1(n823), .A2(n851), .A3(n822), .A4(n821), .Y(n838) );
  AO22X1_LVT U927 ( .A1(n66), .A2(link_addr[16]), .A3(n957), .A4(n890), .Y(
        n824) );
  INVX1_LVT U928 ( .A(n824), .Y(n833) );
  NAND3X0_LVT U929 ( .A1(ex_aluop[0]), .A2(n1127), .A3(opv2[16]), .Y(n825) );
  AND2X1_LVT U930 ( .A1(n825), .A2(n1088), .Y(n827) );
  OR2X1_LVT U931 ( .A1(opv2[16]), .A2(n1127), .Y(n826) );
  AO222X1_LVT U934 ( .A1(n891), .A2(n15), .A3(n829), .A4(n19), .A5(n892), .A6(
        n1083), .Y(n830) );
  NAND2X0_LVT U935 ( .A1(n1086), .A2(n830), .Y(n831) );
  NAND3X0_LVT U936 ( .A1(n833), .A2(n1103), .A3(n831), .Y(n837) );
  INVX1_LVT U937 ( .A(n879), .Y(n848) );
  AO22X1_LVT U938 ( .A1(n1085), .A2(n848), .A3(n1090), .A4(n834), .Y(n836) );
  AO222X1_LVT U940 ( .A1(n926), .A2(n15), .A3(n839), .A4(n19), .A5(n925), .A6(
        n1084), .Y(n841) );
  AO22X1_LVT U941 ( .A1(n1086), .A2(n841), .A3(n957), .A4(n999), .Y(n858) );
  NAND3X0_LVT U942 ( .A1(n1031), .A2(n1133), .A3(opv2[17]), .Y(n842) );
  OA21X1_LVT U943 ( .A1(n1133), .A2(opv2[17]), .A3(n842), .Y(n843) );
  AO22X1_LVT U944 ( .A1(n66), .A2(link_addr[17]), .A3(n1088), .A4(n843), .Y(
        n857) );
  FADDX1_LVT U945 ( .A(opv1[17]), .B(n845), .CI(n844), .CO(n368), .S(n855) );
  NAND2X0_LVT U946 ( .A1(n868), .A2(n846), .Y(n853) );
  NAND4X0_LVT U947 ( .A1(n1031), .A2(n1133), .A3(opv2[17]), .A4(n1087), .Y(
        n852) );
  AOI22X1_LVT U948 ( .A1(n1090), .A2(n849), .A3(n848), .A4(n847), .Y(n850) );
  NAND4X0_LVT U949 ( .A1(n853), .A2(n852), .A3(n851), .A4(n850), .Y(n854) );
  AO21X1_LVT U950 ( .A1(n52), .A2(n855), .A3(n854), .Y(n856) );
  AO222X1_LVT U952 ( .A1(n861), .A2(n15), .A3(n860), .A4(n19), .A5(n961), .A6(
        n1083), .Y(n863) );
  AO22X1_LVT U953 ( .A1(n1086), .A2(n863), .A3(n1090), .A4(n862), .Y(n872) );
  FADDX1_LVT U954 ( .A(opv1[19]), .B(n865), .CI(n864), .CO(n884), .S(n866) );
  AND2X1_LVT U955 ( .A1(n52), .A2(n866), .Y(n871) );
  AO22X1_LVT U956 ( .A1(n957), .A2(n962), .A3(n868), .A4(n867), .Y(n869) );
  AO21X1_LVT U957 ( .A1(n66), .A2(link_addr[19]), .A3(n869), .Y(n870) );
  NOR4X1_LVT U958 ( .A1(n872), .A2(n919), .A3(n871), .A4(n870), .Y(n880) );
  NAND2X0_LVT U959 ( .A1(n1060), .A2(n1062), .Y(n876) );
  NAND3X0_LVT U960 ( .A1(ex_aluop[0]), .A2(n1135), .A3(opv2[19]), .Y(n875) );
  NAND3X0_LVT U961 ( .A1(n1088), .A2(n876), .A3(n875), .Y(n878) );
  NAND4X0_LVT U962 ( .A1(ex_aluop[0]), .A2(n1135), .A3(opv2[19]), .A4(n1087), 
        .Y(n877) );
  NAND3X0_LVT U964 ( .A1(n1031), .A2(n1128), .A3(opv2[20]), .Y(n883) );
  OA21X1_LVT U965 ( .A1(n1128), .A2(opv2[20]), .A3(n883), .Y(n881) );
  AO22X1_LVT U966 ( .A1(n66), .A2(link_addr[20]), .A3(n1088), .A4(n881), .Y(
        n897) );
  INVX1_LVT U967 ( .A(n883), .Y(n888) );
  FADDX1_LVT U968 ( .A(opv1[20]), .B(n885), .CI(n884), .CO(n907), .S(n887) );
  AO222X1_LVT U969 ( .A1(n1087), .A2(n888), .A3(n887), .A4(n52), .A5(n957), 
        .A6(n886), .Y(n896) );
  AO222X1_LVT U970 ( .A1(n892), .A2(n15), .A3(n891), .A4(n19), .A5(n890), .A6(
        n1083), .Y(n894) );
  AO22X1_LVT U971 ( .A1(n1086), .A2(n894), .A3(n1090), .A4(n893), .Y(n895) );
  NOR4X1_LVT U972 ( .A1(n919), .A2(n897), .A3(n896), .A4(n895), .Y(n903) );
  NAND3X0_LVT U973 ( .A1(n899), .A2(n1013), .A3(n1040), .Y(n902) );
  NAND3X0_LVT U974 ( .A1(n987), .A2(n904), .A3(n900), .Y(n901) );
  AND2X1_LVT U976 ( .A1(n987), .A2(n904), .Y(n906) );
  AO22X1_LVT U977 ( .A1(n906), .A2(n986), .A3(n1013), .A4(n905), .Y(n932) );
  FADDX1_LVT U978 ( .A(opv1[21]), .B(n908), .CI(n907), .CO(n383), .S(n916) );
  NAND3X0_LVT U979 ( .A1(ex_aluop[0]), .A2(n1119), .A3(opv2[21]), .Y(n909) );
  INVX1_LVT U980 ( .A(n909), .Y(n914) );
  AND2X1_LVT U981 ( .A1(n909), .A2(n1088), .Y(n911) );
  OR2X1_LVT U982 ( .A1(opv2[21]), .A2(n1119), .Y(n910) );
  AND2X1_LVT U983 ( .A1(n911), .A2(n910), .Y(n912) );
  AO21X1_LVT U984 ( .A1(n66), .A2(link_addr[21]), .A3(n912), .Y(n913) );
  AO21X1_LVT U985 ( .A1(n1087), .A2(n914), .A3(n913), .Y(n915) );
  INVX1_LVT U988 ( .A(n919), .Y(n921) );
  NAND2X0_LVT U989 ( .A1(n957), .A2(n994), .Y(n920) );
  NAND3X0_LVT U990 ( .A1(n1102), .A2(n921), .A3(n920), .Y(n931) );
  AO222X1_LVT U991 ( .A1(n926), .A2(n19), .A3(n925), .A4(n15), .A5(n999), .A6(
        n1083), .Y(n929) );
  AO22X1_LVT U992 ( .A1(n1086), .A2(n929), .A3(n1090), .A4(n927), .Y(n930) );
  AOI22X1_LVT U994 ( .A1(n957), .A2(n934), .A3(n933), .A4(n954), .Y(n953) );
  FADDX1_LVT U995 ( .A(n1124), .B(n936), .CI(n935), .CO(n958), .S(n937) );
  NAND2X0_LVT U996 ( .A1(n52), .A2(n937), .Y(n944) );
  OA221X1_LVT U997 ( .A1(n1124), .A2(n975), .A3(n1071), .A4(n973), .A5(n972), 
        .Y(n941) );
  OA22X1_LVT U998 ( .A1(n941), .A2(n1069), .A3(n939), .A4(n975), .Y(n943) );
  NAND2X0_LVT U999 ( .A1(n66), .A2(link_addr[26]), .Y(n942) );
  AND4X1_LVT U1000 ( .A1(n944), .A2(n943), .A3(n970), .A4(n942), .Y(n952) );
  AOI222X1_LVT U1001 ( .A1(n1084), .A2(n947), .A3(n15), .A4(n946), .A5(n19), 
        .A6(n945), .Y(n948) );
  OA22X1_LVT U1002 ( .A1(n949), .A2(n976), .A3(n948), .A4(n1118), .Y(n951) );
  NAND2X0_LVT U1003 ( .A1(n950), .A2(n987), .Y(n980) );
  AOI22X1_LVT U1005 ( .A1(n957), .A2(n956), .A3(n955), .A4(n954), .Y(n983) );
  FADDX1_LVT U1006 ( .A(n1141), .B(n959), .CI(n958), .CO(n526), .S(n960) );
  NAND2X0_LVT U1007 ( .A1(n52), .A2(n960), .Y(n971) );
  AOI222X1_LVT U1008 ( .A1(n963), .A2(n1084), .A3(n962), .A4(n15), .A5(n961), 
        .A6(n19), .Y(n966) );
  OA22X1_LVT U1009 ( .A1(n966), .A2(n1118), .A3(n964), .A4(n975), .Y(n969) );
  NAND2X0_LVT U1010 ( .A1(n66), .A2(link_addr[27]), .Y(n968) );
  AND4X1_LVT U1011 ( .A1(n971), .A2(n970), .A3(n969), .A4(n968), .Y(n982) );
  OA221X1_LVT U1012 ( .A1(n1141), .A2(n975), .A3(n1070), .A4(n973), .A5(n972), 
        .Y(n979) );
  OA22X1_LVT U1013 ( .A1(n979), .A2(n1068), .A3(n977), .A4(n976), .Y(n981) );
  AOI22X1_LVT U1015 ( .A1(n987), .A2(n986), .A3(n985), .A4(n984), .Y(n1028) );
  FADDX1_LVT U1016 ( .A(opv1[29]), .B(n989), .CI(n988), .CO(n559), .S(n1023)
         );
  NAND3X0_LVT U1017 ( .A1(ex_aluop[0]), .A2(opv1[29]), .A3(opv2[29]), .Y(n991)
         );
  AND2X1_LVT U1018 ( .A1(n991), .A2(n1088), .Y(n993) );
  OR2X1_LVT U1019 ( .A1(opv2[29]), .A2(opv1[29]), .Y(n992) );
  AND2X1_LVT U1020 ( .A1(n993), .A2(n992), .Y(n1020) );
  AO22X1_LVT U1021 ( .A1(n1084), .A2(n996), .A3(n15), .A4(n994), .Y(n998) );
  INVX1_LVT U1022 ( .A(n998), .Y(n1011) );
  AO22X1_LVT U1023 ( .A1(n1001), .A2(opv1[29]), .A3(n19), .A4(n999), .Y(n1002)
         );
  INVX1_LVT U1024 ( .A(n1002), .Y(n1010) );
  NAND2X0_LVT U1025 ( .A1(n1140), .A2(n16), .Y(n1005) );
  NAND3X0_LVT U1026 ( .A1(n1006), .A2(n1005), .A3(n1004), .Y(n1007) );
  NAND2X0_LVT U1027 ( .A1(n28), .A2(n1007), .Y(n1009) );
  NAND3X0_LVT U1028 ( .A1(n1011), .A2(n1010), .A3(n1009), .Y(n1014) );
  AO22X1_LVT U1029 ( .A1(n1086), .A2(n1014), .A3(n1013), .A4(n1012), .Y(n1016)
         );
  AO21X1_LVT U1030 ( .A1(n66), .A2(link_addr[29]), .A3(n1016), .Y(n1018) );
  OR3X1_LVT U1031 ( .A1(n1020), .A2(n1019), .A3(n1018), .Y(n1021) );
  NAND4X0_LVT U1034 ( .A1(ex_aluop[0]), .A2(opv1[29]), .A3(opv2[29]), .A4(
        n1087), .Y(n1026) );
  AO21X2_LVT U754 ( .A1(n602), .A2(n52), .A3(n601), .Y(reg_wdata[31]) );
  NAND4X0_LVT U1014 ( .A1(n983), .A2(n982), .A3(n981), .A4(n980), .Y(
        reg_wdata[27]) );
  AO21X2_LVT U724 ( .A1(n558), .A2(n52), .A3(n557), .Y(reg_wdata[28]) );
  NAND4X0_LVT U1004 ( .A1(n953), .A2(n952), .A3(n951), .A4(n980), .Y(
        reg_wdata[26]) );
  AO21X2_LVT U695 ( .A1(n52), .A2(n525), .A3(n524), .Y(reg_wdata[25]) );
  AO21X2_LVT U673 ( .A1(n52), .A2(n487), .A3(n486), .Y(reg_wdata[24]) );
  AO21X2_LVT U648 ( .A1(n52), .A2(n442), .A3(n441), .Y(reg_wdata[23]) );
  NAND4X0_LVT U963 ( .A1(n880), .A2(n879), .A3(n878), .A4(n877), .Y(
        reg_wdata[19]) );
  NAND4X0_LVT U612 ( .A1(n382), .A2(n381), .A3(n879), .A4(n380), .Y(
        reg_wdata[18]) );
  NAND4X0_LVT U921 ( .A1(n817), .A2(n816), .A3(n815), .A4(n851), .Y(
        reg_wdata[15]) );
  NAND4X0_LVT U494 ( .A1(n252), .A2(n251), .A3(n250), .A4(n249), .Y(
        reg_wdata[0]) );
  NAND2X2_LVT U873 ( .A1(n741), .A2(n740), .Y(reg_wdata[11]) );
  NAND4X0_LVT U546 ( .A1(n303), .A2(n302), .A3(n301), .A4(n1099), .Y(
        reg_wdata[2]) );
  NOR2X4_LVT U16 ( .A1(n6), .A2(n5), .Y(n52) );
  NAND2X0_LVT U162 ( .A1(aluop[1]), .A2(n65), .Y(n975) );
  NAND4X0_LVT U79 ( .A1(n1031), .A2(n430), .A3(n1034), .A4(n1042), .Y(n965) );
  AND2X4_LVT U68 ( .A1(n1040), .A2(n1038), .Y(n28) );
  AND2X4_LVT U84 ( .A1(N287), .A2(n1036), .Y(n16) );
  AND2X4_LVT U97 ( .A1(opv2[3]), .A2(n1038), .Y(n15) );
  AND3X4_LVT U181 ( .A1(alusel[2]), .A2(alusel[1]), .A3(n48), .Y(n66) );
  AND4X2_LVT U52 ( .A1(aluop[2]), .A2(alusel[1]), .A3(n8), .A4(n48), .Y(n430)
         );
  AND2X4_LVT U110 ( .A1(opv2[3]), .A2(opv2[2]), .Y(n19) );
  AND4X4_LVT U347 ( .A1(alusel[2]), .A2(alusel[0]), .A3(alusel[1]), .A4(n1030), 
        .Y(n130) );
  INVX1_LVT U3 ( .A(rst), .Y(n1030) );
  NBUFFX4_LVT U4 ( .A(aluop[0]), .Y(n1031) );
  NBUFFX4_LVT U5 ( .A(aluop[0]), .Y(ex_aluop[0]) );
  INVX1_LVT U11 ( .A(ex_aluop[0]), .Y(n1033) );
  INVX1_LVT U12 ( .A(aluop[1]), .Y(n1034) );
  INVX2_LVT U13 ( .A(N287), .Y(n1035) );
  INVX1_LVT U17 ( .A(opv2[1]), .Y(n1036) );
  INVX1_LVT U18 ( .A(opv1[0]), .Y(n1037) );
  INVX1_LVT U53 ( .A(opv1[1]), .Y(n1039) );
  INVX2_LVT U54 ( .A(opv2[3]), .Y(n1040) );
  INVX1_LVT U55 ( .A(n1122), .Y(n1041) );
  INVX2_LVT U57 ( .A(opv2[4]), .Y(n1042) );
  INVX1_LVT U58 ( .A(n1142), .Y(n1043) );
  INVX1_LVT U59 ( .A(n1114), .Y(n1044) );
  INVX1_LVT U60 ( .A(n1137), .Y(n1045) );
  INVX1_LVT U61 ( .A(n1125), .Y(n1046) );
  INVX1_LVT U64 ( .A(n1126), .Y(n1047) );
  INVX1_LVT U69 ( .A(n1129), .Y(n1048) );
  INVX1_LVT U73 ( .A(n1123), .Y(n1049) );
  INVX1_LVT U78 ( .A(opv2[11]), .Y(n1050) );
  INVX1_LVT U80 ( .A(n1136), .Y(n1051) );
  INVX1_LVT U82 ( .A(n1132), .Y(n1052) );
  INVX1_LVT U83 ( .A(n1116), .Y(n1053) );
  INVX1_LVT U85 ( .A(n1134), .Y(n1054) );
  INVX1_LVT U88 ( .A(opv2[15]), .Y(n1055) );
  INVX1_LVT U89 ( .A(n1117), .Y(n1056) );
  INVX1_LVT U93 ( .A(n1120), .Y(n1057) );
  INVX1_LVT U94 ( .A(n1127), .Y(n1058) );
  INVX1_LVT U98 ( .A(n1133), .Y(n1059) );
  INVX1_LVT U99 ( .A(opv2[19]), .Y(n1060) );
  INVX1_LVT U100 ( .A(n1130), .Y(n1061) );
  INVX1_LVT U102 ( .A(n1135), .Y(n1062) );
  INVX1_LVT U104 ( .A(n1128), .Y(n1063) );
  INVX1_LVT U111 ( .A(opv2[22]), .Y(n1064) );
  INVX1_LVT U112 ( .A(n1119), .Y(n1065) );
  INVX1_LVT U126 ( .A(opv1[23]), .Y(n1066) );
  INVX1_LVT U136 ( .A(opv1[22]), .Y(n1067) );
  INVX1_LVT U142 ( .A(opv2[27]), .Y(n1068) );
  INVX1_LVT U143 ( .A(opv2[26]), .Y(n1069) );
  INVX1_LVT U144 ( .A(opv1[27]), .Y(n1070) );
  INVX1_LVT U163 ( .A(opv1[26]), .Y(n1071) );
  INVX1_LVT U164 ( .A(opv1[24]), .Y(n1072) );
  INVX1_LVT U165 ( .A(opv1[25]), .Y(n1073) );
  INVX1_LVT U166 ( .A(n1143), .Y(n1074) );
  INVX1_LVT U182 ( .A(opv1[28]), .Y(n1075) );
  INVX1_LVT U185 ( .A(opv2[28]), .Y(n1076) );
  INVX1_LVT U191 ( .A(opv2[29]), .Y(n1077) );
  INVX1_LVT U199 ( .A(opv2[30]), .Y(n1078) );
  INVX1_LVT U206 ( .A(opv2[31]), .Y(n1079) );
  INVX4_LVT U208 ( .A(n86), .Y(n1080) );
  INVX1_LVT U209 ( .A(n430), .Y(n1081) );
  INVX4_LVT U229 ( .A(n29), .Y(n1082) );
  NBUFFX4_LVT U235 ( .A(n13), .Y(n1083) );
  NBUFFX4_LVT U250 ( .A(n13), .Y(n1084) );
  INVX4_LVT U256 ( .A(n176), .Y(n1085) );
  INVX4_LVT U346 ( .A(n965), .Y(n1086) );
  INVX4_LVT U348 ( .A(n798), .Y(n1087) );
  INVX4_LVT U349 ( .A(n975), .Y(n1088) );
  INVX1_LVT U385 ( .A(n1139), .Y(n1089) );
  INVX2_LVT U388 ( .A(n812), .Y(n1090) );
  OR3X2_LVT U835 ( .A1(n690), .A2(n689), .A3(n688), .Y(reg_wdata[4]) );
  OR3X2_LVT U888 ( .A1(n763), .A2(n762), .A3(n761), .Y(reg_wdata[12]) );
  OR3X2_LVT U993 ( .A1(n932), .A2(n931), .A3(n930), .Y(reg_wdata[21]) );
  AO21X2_LVT U520 ( .A1(n52), .A2(n278), .A3(n277), .Y(reg_wdata[1]) );
  OR3X2_LVT U850 ( .A1(n707), .A2(n706), .A3(n705), .Y(reg_wdata[5]) );
  OR3X2_LVT U951 ( .A1(n858), .A2(n857), .A3(n856), .Y(reg_wdata[17]) );
  OR3X2_LVT U906 ( .A1(n789), .A2(n788), .A3(n787), .Y(reg_wdata[13]) );
  OR3X2_LVT U939 ( .A1(n838), .A2(n837), .A3(n836), .Y(reg_wdata[16]) );
  OR3X2_LVT U861 ( .A1(n723), .A2(n722), .A3(n721), .Y(reg_wdata[8]) );
  AO21X2_LVT U562 ( .A1(n52), .A2(n324), .A3(n323), .Y(reg_wdata[3]) );
  AO21X2_LVT U628 ( .A1(n52), .A2(n405), .A3(n404), .Y(reg_wdata[22]) );
  AO21X2_LVT U580 ( .A1(n52), .A2(n343), .A3(n342), .Y(reg_wdata[6]) );
  AO21X2_LVT U599 ( .A1(n52), .A2(n367), .A3(n366), .Y(reg_wdata[14]) );
  INVX4_LVT U43 ( .A(opv2[2]), .Y(n1038) );
  NAND3X2_LVT U344 ( .A1(n1101), .A2(n1100), .A3(n126), .Y(reg_wdata[7]) );
  NAND3X2_LVT U975 ( .A1(n903), .A2(n902), .A3(n901), .Y(reg_wdata[20]) );
  NAND3X2_LVT U288 ( .A1(n1106), .A2(n1107), .A3(n101), .Y(reg_wdata[9]) );
  AND2X4_LVT U10 ( .A1(n1031), .A2(aluop[1]), .Y(n2) );
  INVX2_LVT U63 ( .A(n88), .Y(n1001) );
  NAND3X2_LVT U228 ( .A1(n1108), .A2(n77), .A3(n76), .Y(reg_wdata[10]) );
  NAND3X2_LVT U1035 ( .A1(n1028), .A2(n1109), .A3(n1026), .Y(reg_wdata[29]) );
  NBUFFX4_LVT U158 ( .A(opv1[4]), .Y(n1114) );
  NBUFFX4_LVT U159 ( .A(opv1[2]), .Y(n1122) );
  NBUFFX4_LVT U179 ( .A(opv1[3]), .Y(n1142) );
  NBUFFX4_LVT U180 ( .A(opv1[14]), .Y(n1117) );
  NBUFFX4_LVT U214 ( .A(opv1[13]), .Y(n1134) );
  NBUFFX4_LVT U215 ( .A(opv1[9]), .Y(n1123) );
  NBUFFX4_LVT U275 ( .A(opv1[5]), .Y(n1137) );
  NBUFFX4_LVT U276 ( .A(opv1[10]), .Y(n1136) );
  NBUFFX4_LVT U278 ( .A(opv1[12]), .Y(n1116) );
  NBUFFX4_LVT U279 ( .A(opv1[6]), .Y(n1125) );
  NBUFFX4_LVT U299 ( .A(opv1[15]), .Y(n1120) );
  NBUFFX4_LVT U300 ( .A(opv1[8]), .Y(n1129) );
  NBUFFX4_LVT U312 ( .A(opv1[7]), .Y(n1126) );
  NBUFFX4_LVT U313 ( .A(opv1[11]), .Y(n1132) );
  NBUFFX4_LVT U325 ( .A(opv1[18]), .Y(n1130) );
  NBUFFX4_LVT U326 ( .A(opv1[21]), .Y(n1119) );
  NBUFFX4_LVT U389 ( .A(opv1[17]), .Y(n1133) );
  NBUFFX4_LVT U390 ( .A(opv1[20]), .Y(n1128) );
  NBUFFX4_LVT U393 ( .A(opv1[16]), .Y(n1127) );
  NBUFFX4_LVT U394 ( .A(opv1[19]), .Y(n1135) );
  NBUFFX4_LVT U397 ( .A(opv1[22]), .Y(n1113) );
  NBUFFX4_LVT U398 ( .A(opv1[24]), .Y(n1115) );
  NBUFFX4_LVT U399 ( .A(opv1[23]), .Y(n1112) );
  NBUFFX4_LVT U402 ( .A(opv1[25]), .Y(n1121) );
  NBUFFX4_LVT U404 ( .A(opv1[30]), .Y(n1131) );
  NBUFFX4_LVT U408 ( .A(opv1[26]), .Y(n1124) );
  NBUFFX4_LVT U409 ( .A(opv1[27]), .Y(n1141) );
  NBUFFX4_LVT U410 ( .A(opv1[28]), .Y(n1140) );
  NAND2X0_LVT U413 ( .A1(n332), .A2(n331), .Y(n1091) );
  NAND2X0_LVT U415 ( .A1(n286), .A2(n285), .Y(n1092) );
  NAND2X0_LVT U419 ( .A1(n268), .A2(n267), .Y(n1093) );
  AOI22X1_LVT U420 ( .A1(n66), .A2(link_addr[2]), .A3(n957), .A4(n373), .Y(
        n1094) );
  NAND2X0_LVT U421 ( .A1(n109), .A2(n108), .Y(n1095) );
  NAND2X0_LVT U424 ( .A1(n356), .A2(n355), .Y(n1096) );
  AND3X1_LVT U426 ( .A1(n511), .A2(n510), .A3(n970), .Y(n1097) );
  AOI22X1_LVT U430 ( .A1(n1086), .A2(n505), .A3(n1013), .A4(n504), .Y(n1098)
         );
  AND3X1_LVT U431 ( .A1(n1094), .A2(n1092), .A3(n296), .Y(n1099) );
  AND4X1_LVT U432 ( .A1(n123), .A2(n122), .A3(n121), .A4(n120), .Y(n1100) );
  AND3X1_LVT U440 ( .A1(n113), .A2(n1095), .A3(n111), .Y(n1101) );
  AOI21X1_LVT U443 ( .A1(n52), .A2(n916), .A3(n915), .Y(n1102) );
  NAND2X0_LVT U445 ( .A1(n827), .A2(n826), .Y(n1103) );
  AOI21X1_LVT U451 ( .A1(n52), .A2(n774), .A3(n773), .Y(n1104) );
  AOI21X1_LVT U453 ( .A1(n52), .A2(n751), .A3(n750), .Y(n1105) );
  AOI222X1_LVT U454 ( .A1(n95), .A2(n430), .A3(n52), .A4(n94), .A5(n93), .A6(
        n1087), .Y(n1106) );
  AOI22X1_LVT U457 ( .A1(n66), .A2(link_addr[9]), .A3(n1088), .A4(n98), .Y(
        n1107) );
  AOI21X1_LVT U470 ( .A1(n52), .A2(n74), .A3(n73), .Y(n1108) );
  AOI21X1_LVT U472 ( .A1(n1023), .A2(n52), .A3(n1021), .Y(n1109) );
  AOI221X1_LVT U478 ( .A1(n1088), .A2(n46), .A3(n1088), .A4(n230), .A5(n45), 
        .Y(n1110) );
  AOI21X1_LVT U484 ( .A1(n52), .A2(n35), .A3(n34), .Y(n1111) );
  NBUFFX4_LVT U513 ( .A(n130), .Y(n1144) );
  NBUFFX4_LVT U514 ( .A(opv2[9]), .Y(rt_data[9]) );
  NBUFFX4_LVT U527 ( .A(n965), .Y(n1118) );
  NBUFFX4_LVT U528 ( .A(n2), .Y(n1139) );
  NBUFFX4_LVT U531 ( .A(opv1[31]), .Y(n1143) );
endmodule


module pipe_ex_mem ( clk, rst, ex_reg_waddr, ex_we, ex_reg_wdata, stall, 
        ex_mem_addr, ex_aluop, ex_rt_data, mem_reg_waddr, mem_we, 
        mem_reg_wdata, mem_mem_addr, mem_aluop, mem_rt_data );
  input [4:0] ex_reg_waddr;
  input [31:0] ex_reg_wdata;
  input [5:0] stall;
  input [31:0] ex_mem_addr;
  input [7:0] ex_aluop;
  input [31:0] ex_rt_data;
  output [4:0] mem_reg_waddr;
  output [31:0] mem_reg_wdata;
  output [31:0] mem_mem_addr;
  output [7:0] mem_aluop;
  output [31:0] mem_rt_data;
  input clk, rst, ex_we;
  output mem_we;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n2, n3, n135,
         n136, n137, n138, n139, n140, n141, n143;

  DFFX1_LVT \mem_rt_data_reg[31]  ( .D(n73), .CLK(clk), .Q(mem_rt_data[31]) );
  DFFX1_LVT \mem_rt_data_reg[30]  ( .D(n72), .CLK(clk), .Q(mem_rt_data[30]) );
  DFFX1_LVT \mem_rt_data_reg[29]  ( .D(n71), .CLK(clk), .Q(mem_rt_data[29]) );
  DFFX1_LVT \mem_rt_data_reg[28]  ( .D(n70), .CLK(clk), .Q(mem_rt_data[28]) );
  DFFX1_LVT \mem_rt_data_reg[27]  ( .D(n69), .CLK(clk), .Q(mem_rt_data[27]) );
  DFFX1_LVT \mem_rt_data_reg[26]  ( .D(n68), .CLK(clk), .Q(mem_rt_data[26]) );
  DFFX1_LVT \mem_rt_data_reg[25]  ( .D(n67), .CLK(clk), .Q(mem_rt_data[25]) );
  DFFX1_LVT \mem_rt_data_reg[24]  ( .D(n66), .CLK(clk), .Q(mem_rt_data[24]) );
  DFFX1_LVT \mem_rt_data_reg[23]  ( .D(n65), .CLK(clk), .Q(mem_rt_data[23]) );
  DFFX1_LVT \mem_rt_data_reg[22]  ( .D(n64), .CLK(clk), .Q(mem_rt_data[22]) );
  DFFX1_LVT \mem_rt_data_reg[21]  ( .D(n63), .CLK(clk), .Q(mem_rt_data[21]) );
  DFFX1_LVT \mem_rt_data_reg[20]  ( .D(n62), .CLK(clk), .Q(mem_rt_data[20]) );
  DFFX1_LVT \mem_rt_data_reg[19]  ( .D(n61), .CLK(clk), .Q(mem_rt_data[19]) );
  DFFX1_LVT \mem_rt_data_reg[18]  ( .D(n60), .CLK(clk), .Q(mem_rt_data[18]) );
  DFFX1_LVT \mem_rt_data_reg[17]  ( .D(n59), .CLK(clk), .Q(mem_rt_data[17]) );
  DFFX1_LVT \mem_rt_data_reg[16]  ( .D(n58), .CLK(clk), .Q(mem_rt_data[16]) );
  DFFX1_LVT \mem_reg_waddr_reg[4]  ( .D(n41), .CLK(clk), .Q(mem_reg_waddr[4])
         );
  DFFX1_LVT \mem_reg_waddr_reg[3]  ( .D(n40), .CLK(clk), .Q(mem_reg_waddr[3])
         );
  DFFX1_LVT \mem_reg_waddr_reg[2]  ( .D(n39), .CLK(clk), .Q(mem_reg_waddr[2])
         );
  DFFX1_LVT \mem_reg_waddr_reg[1]  ( .D(n38), .CLK(clk), .Q(mem_reg_waddr[1])
         );
  DFFX1_LVT \mem_reg_waddr_reg[0]  ( .D(n37), .CLK(clk), .Q(mem_reg_waddr[0])
         );
  DFFX1_LVT mem_we_reg ( .D(n36), .CLK(clk), .Q(mem_we) );
  DFFX1_LVT \mem_reg_wdata_reg[14]  ( .D(n18), .CLK(clk), .Q(mem_reg_wdata[14]) );
  DFFX1_LVT \mem_reg_wdata_reg[13]  ( .D(n17), .CLK(clk), .Q(mem_reg_wdata[13]) );
  DFFX1_LVT \mem_reg_wdata_reg[12]  ( .D(n16), .CLK(clk), .Q(mem_reg_wdata[12]) );
  DFFX1_LVT \mem_reg_wdata_reg[11]  ( .D(n15), .CLK(clk), .Q(mem_reg_wdata[11]) );
  DFFX1_LVT \mem_reg_wdata_reg[10]  ( .D(n14), .CLK(clk), .Q(mem_reg_wdata[10]) );
  DFFX1_LVT \mem_reg_wdata_reg[9]  ( .D(n13), .CLK(clk), .Q(mem_reg_wdata[9])
         );
  DFFX1_LVT \mem_reg_wdata_reg[8]  ( .D(n12), .CLK(clk), .Q(mem_reg_wdata[8])
         );
  DFFX1_LVT \mem_reg_wdata_reg[7]  ( .D(n11), .CLK(clk), .Q(mem_reg_wdata[7])
         );
  DFFX1_LVT \mem_reg_wdata_reg[31]  ( .D(n35), .CLK(clk), .Q(mem_reg_wdata[31]) );
  DFFX1_LVT \mem_reg_wdata_reg[30]  ( .D(n34), .CLK(clk), .Q(mem_reg_wdata[30]) );
  DFFX1_LVT \mem_reg_wdata_reg[29]  ( .D(n33), .CLK(clk), .Q(mem_reg_wdata[29]) );
  DFFX1_LVT \mem_reg_wdata_reg[28]  ( .D(n32), .CLK(clk), .Q(mem_reg_wdata[28]) );
  DFFX1_LVT \mem_reg_wdata_reg[27]  ( .D(n31), .CLK(clk), .Q(mem_reg_wdata[27]) );
  DFFX1_LVT \mem_reg_wdata_reg[26]  ( .D(n30), .CLK(clk), .Q(mem_reg_wdata[26]) );
  DFFX1_LVT \mem_reg_wdata_reg[25]  ( .D(n29), .CLK(clk), .Q(mem_reg_wdata[25]) );
  DFFX1_LVT \mem_reg_wdata_reg[24]  ( .D(n28), .CLK(clk), .Q(mem_reg_wdata[24]) );
  DFFX1_LVT \mem_reg_wdata_reg[23]  ( .D(n27), .CLK(clk), .Q(mem_reg_wdata[23]) );
  DFFX1_LVT \mem_reg_wdata_reg[22]  ( .D(n26), .CLK(clk), .Q(mem_reg_wdata[22]) );
  DFFX1_LVT \mem_reg_wdata_reg[21]  ( .D(n25), .CLK(clk), .Q(mem_reg_wdata[21]) );
  DFFX1_LVT \mem_reg_wdata_reg[20]  ( .D(n24), .CLK(clk), .Q(mem_reg_wdata[20]) );
  DFFX1_LVT \mem_reg_wdata_reg[19]  ( .D(n23), .CLK(clk), .Q(mem_reg_wdata[19]) );
  DFFX1_LVT \mem_reg_wdata_reg[18]  ( .D(n22), .CLK(clk), .Q(mem_reg_wdata[18]) );
  DFFX1_LVT \mem_reg_wdata_reg[17]  ( .D(n21), .CLK(clk), .Q(mem_reg_wdata[17]) );
  DFFX1_LVT \mem_reg_wdata_reg[16]  ( .D(n20), .CLK(clk), .Q(mem_reg_wdata[16]) );
  DFFX1_LVT \mem_reg_wdata_reg[15]  ( .D(n19), .CLK(clk), .Q(mem_reg_wdata[15]) );
  DFFX1_LVT \mem_mem_addr_reg[31]  ( .D(n113), .CLK(clk), .Q(mem_mem_addr[31])
         );
  DFFX1_LVT \mem_mem_addr_reg[30]  ( .D(n112), .CLK(clk), .Q(mem_mem_addr[30])
         );
  DFFX1_LVT \mem_mem_addr_reg[29]  ( .D(n111), .CLK(clk), .Q(mem_mem_addr[29])
         );
  DFFX1_LVT \mem_mem_addr_reg[28]  ( .D(n110), .CLK(clk), .Q(mem_mem_addr[28])
         );
  DFFX1_LVT \mem_mem_addr_reg[27]  ( .D(n109), .CLK(clk), .Q(mem_mem_addr[27])
         );
  DFFX1_LVT \mem_mem_addr_reg[26]  ( .D(n108), .CLK(clk), .Q(mem_mem_addr[26])
         );
  DFFX1_LVT \mem_mem_addr_reg[25]  ( .D(n107), .CLK(clk), .Q(mem_mem_addr[25])
         );
  DFFX1_LVT \mem_mem_addr_reg[24]  ( .D(n106), .CLK(clk), .Q(mem_mem_addr[24])
         );
  DFFX1_LVT \mem_mem_addr_reg[23]  ( .D(n105), .CLK(clk), .Q(mem_mem_addr[23])
         );
  DFFX1_LVT \mem_mem_addr_reg[22]  ( .D(n104), .CLK(clk), .Q(mem_mem_addr[22])
         );
  DFFX1_LVT \mem_mem_addr_reg[21]  ( .D(n103), .CLK(clk), .Q(mem_mem_addr[21])
         );
  DFFX1_LVT \mem_mem_addr_reg[20]  ( .D(n102), .CLK(clk), .Q(mem_mem_addr[20])
         );
  DFFX1_LVT \mem_mem_addr_reg[19]  ( .D(n101), .CLK(clk), .Q(mem_mem_addr[19])
         );
  DFFX1_LVT \mem_mem_addr_reg[18]  ( .D(n100), .CLK(clk), .Q(mem_mem_addr[18])
         );
  DFFX1_LVT \mem_mem_addr_reg[17]  ( .D(n99), .CLK(clk), .Q(mem_mem_addr[17])
         );
  DFFX1_LVT \mem_mem_addr_reg[16]  ( .D(n98), .CLK(clk), .Q(mem_mem_addr[16])
         );
  DFFX1_LVT \mem_mem_addr_reg[15]  ( .D(n97), .CLK(clk), .Q(mem_mem_addr[15])
         );
  DFFX1_LVT \mem_mem_addr_reg[14]  ( .D(n96), .CLK(clk), .Q(mem_mem_addr[14])
         );
  DFFX1_LVT \mem_mem_addr_reg[13]  ( .D(n95), .CLK(clk), .Q(mem_mem_addr[13])
         );
  DFFX1_LVT \mem_mem_addr_reg[12]  ( .D(n94), .CLK(clk), .Q(mem_mem_addr[12])
         );
  DFFX1_LVT \mem_mem_addr_reg[11]  ( .D(n93), .CLK(clk), .Q(mem_mem_addr[11])
         );
  DFFX1_LVT \mem_mem_addr_reg[10]  ( .D(n92), .CLK(clk), .Q(mem_mem_addr[10])
         );
  DFFX1_LVT \mem_mem_addr_reg[9]  ( .D(n91), .CLK(clk), .Q(mem_mem_addr[9]) );
  DFFX1_LVT \mem_mem_addr_reg[8]  ( .D(n90), .CLK(clk), .Q(mem_mem_addr[8]) );
  DFFX1_LVT \mem_mem_addr_reg[7]  ( .D(n89), .CLK(clk), .Q(mem_mem_addr[7]) );
  DFFX1_LVT \mem_mem_addr_reg[6]  ( .D(n88), .CLK(clk), .Q(mem_mem_addr[6]) );
  DFFX1_LVT \mem_mem_addr_reg[5]  ( .D(n87), .CLK(clk), .Q(mem_mem_addr[5]) );
  DFFX1_LVT \mem_mem_addr_reg[4]  ( .D(n86), .CLK(clk), .Q(mem_mem_addr[4]) );
  DFFX1_LVT \mem_mem_addr_reg[3]  ( .D(n85), .CLK(clk), .Q(mem_mem_addr[3]) );
  DFFX1_LVT \mem_mem_addr_reg[2]  ( .D(n84), .CLK(clk), .Q(mem_mem_addr[2]) );
  DFFX1_LVT \mem_rt_data_reg[15]  ( .D(n57), .CLK(clk), .Q(mem_rt_data[15]) );
  DFFX1_LVT \mem_rt_data_reg[14]  ( .D(n56), .CLK(clk), .Q(mem_rt_data[14]) );
  DFFX1_LVT \mem_rt_data_reg[13]  ( .D(n55), .CLK(clk), .Q(mem_rt_data[13]) );
  DFFX1_LVT \mem_rt_data_reg[12]  ( .D(n54), .CLK(clk), .Q(mem_rt_data[12]) );
  DFFX1_LVT \mem_rt_data_reg[11]  ( .D(n53), .CLK(clk), .Q(mem_rt_data[11]) );
  DFFX1_LVT \mem_rt_data_reg[10]  ( .D(n52), .CLK(clk), .Q(mem_rt_data[10]) );
  DFFX1_LVT \mem_rt_data_reg[9]  ( .D(n51), .CLK(clk), .Q(mem_rt_data[9]) );
  DFFX1_LVT \mem_rt_data_reg[8]  ( .D(n50), .CLK(clk), .Q(mem_rt_data[8]) );
  DFFX1_LVT \mem_reg_wdata_reg[0]  ( .D(n4), .CLK(clk), .Q(mem_reg_wdata[0])
         );
  DFFX1_LVT \mem_reg_wdata_reg[6]  ( .D(n10), .CLK(clk), .Q(mem_reg_wdata[6])
         );
  DFFX1_LVT \mem_reg_wdata_reg[5]  ( .D(n9), .CLK(clk), .Q(mem_reg_wdata[5])
         );
  DFFX1_LVT \mem_reg_wdata_reg[4]  ( .D(n8), .CLK(clk), .Q(mem_reg_wdata[4])
         );
  DFFX1_LVT \mem_reg_wdata_reg[3]  ( .D(n7), .CLK(clk), .Q(mem_reg_wdata[3])
         );
  DFFX1_LVT \mem_reg_wdata_reg[2]  ( .D(n6), .CLK(clk), .Q(mem_reg_wdata[2])
         );
  DFFX1_LVT \mem_reg_wdata_reg[1]  ( .D(n5), .CLK(clk), .Q(mem_reg_wdata[1])
         );
  DFFX1_LVT \mem_rt_data_reg[7]  ( .D(n49), .CLK(clk), .Q(mem_rt_data[7]) );
  DFFX1_LVT \mem_rt_data_reg[6]  ( .D(n48), .CLK(clk), .Q(mem_rt_data[6]) );
  DFFX1_LVT \mem_rt_data_reg[5]  ( .D(n47), .CLK(clk), .Q(mem_rt_data[5]) );
  DFFX1_LVT \mem_rt_data_reg[0]  ( .D(n42), .CLK(clk), .Q(mem_rt_data[0]) );
  DFFX1_LVT \mem_mem_addr_reg[0]  ( .D(n82), .CLK(clk), .Q(mem_mem_addr[0]) );
  DFFX1_LVT \mem_aluop_reg[4]  ( .D(n78), .CLK(clk), .Q(mem_aluop[4]) );
  DFFX1_LVT \mem_aluop_reg[2]  ( .D(n76), .CLK(clk), .Q(mem_aluop[2]) );
  DFFX1_LVT \mem_aluop_reg[3]  ( .D(n77), .CLK(clk), .Q(mem_aluop[3]) );
  AO22X1_LVT U12 ( .A1(n137), .A2(mem_mem_addr[31]), .A3(n141), .A4(
        ex_mem_addr[31]), .Y(n113) );
  AO22X1_LVT U13 ( .A1(n137), .A2(mem_mem_addr[30]), .A3(n141), .A4(
        ex_mem_addr[30]), .Y(n112) );
  AO22X1_LVT U14 ( .A1(n137), .A2(mem_mem_addr[29]), .A3(n141), .A4(
        ex_mem_addr[29]), .Y(n111) );
  AO22X1_LVT U15 ( .A1(n137), .A2(mem_mem_addr[28]), .A3(n141), .A4(
        ex_mem_addr[28]), .Y(n110) );
  AO22X1_LVT U16 ( .A1(n137), .A2(mem_mem_addr[27]), .A3(n141), .A4(
        ex_mem_addr[27]), .Y(n109) );
  AO22X1_LVT U17 ( .A1(n137), .A2(mem_mem_addr[26]), .A3(n141), .A4(
        ex_mem_addr[26]), .Y(n108) );
  AO22X1_LVT U18 ( .A1(n137), .A2(mem_mem_addr[25]), .A3(n141), .A4(
        ex_mem_addr[25]), .Y(n107) );
  AO22X1_LVT U19 ( .A1(n137), .A2(mem_mem_addr[24]), .A3(n141), .A4(
        ex_mem_addr[24]), .Y(n106) );
  AO22X1_LVT U20 ( .A1(n137), .A2(mem_mem_addr[23]), .A3(n141), .A4(
        ex_mem_addr[23]), .Y(n105) );
  AO22X1_LVT U21 ( .A1(n137), .A2(mem_mem_addr[22]), .A3(n141), .A4(
        ex_mem_addr[22]), .Y(n104) );
  AO22X1_LVT U22 ( .A1(n137), .A2(mem_mem_addr[21]), .A3(n141), .A4(
        ex_mem_addr[21]), .Y(n103) );
  AO22X1_LVT U23 ( .A1(n137), .A2(mem_mem_addr[20]), .A3(n141), .A4(
        ex_mem_addr[20]), .Y(n102) );
  AO22X1_LVT U24 ( .A1(n137), .A2(mem_mem_addr[19]), .A3(n141), .A4(
        ex_mem_addr[19]), .Y(n101) );
  AO22X1_LVT U25 ( .A1(n137), .A2(mem_mem_addr[18]), .A3(n141), .A4(
        ex_mem_addr[18]), .Y(n100) );
  AO22X1_LVT U26 ( .A1(n137), .A2(mem_mem_addr[17]), .A3(n141), .A4(
        ex_mem_addr[17]), .Y(n99) );
  AO22X1_LVT U29 ( .A1(n137), .A2(mem_mem_addr[16]), .A3(n141), .A4(
        ex_mem_addr[16]), .Y(n98) );
  AO22X1_LVT U30 ( .A1(n137), .A2(mem_mem_addr[15]), .A3(n141), .A4(
        ex_mem_addr[15]), .Y(n97) );
  AO22X1_LVT U31 ( .A1(n137), .A2(mem_mem_addr[14]), .A3(n141), .A4(
        ex_mem_addr[14]), .Y(n96) );
  AO22X1_LVT U32 ( .A1(n137), .A2(mem_mem_addr[13]), .A3(n141), .A4(
        ex_mem_addr[13]), .Y(n95) );
  AO22X1_LVT U33 ( .A1(n137), .A2(mem_mem_addr[12]), .A3(n141), .A4(
        ex_mem_addr[12]), .Y(n94) );
  AO22X1_LVT U34 ( .A1(n137), .A2(mem_mem_addr[11]), .A3(n141), .A4(
        ex_mem_addr[11]), .Y(n93) );
  AO22X1_LVT U35 ( .A1(n137), .A2(mem_mem_addr[10]), .A3(n141), .A4(
        ex_mem_addr[10]), .Y(n92) );
  AO22X1_LVT U36 ( .A1(n137), .A2(mem_mem_addr[9]), .A3(n141), .A4(
        ex_mem_addr[9]), .Y(n91) );
  AO22X1_LVT U37 ( .A1(n137), .A2(mem_mem_addr[8]), .A3(n141), .A4(
        ex_mem_addr[8]), .Y(n90) );
  AO22X1_LVT U38 ( .A1(n137), .A2(mem_mem_addr[7]), .A3(n141), .A4(
        ex_mem_addr[7]), .Y(n89) );
  AO22X1_LVT U39 ( .A1(n137), .A2(mem_mem_addr[6]), .A3(n141), .A4(
        ex_mem_addr[6]), .Y(n88) );
  AO22X1_LVT U40 ( .A1(n137), .A2(mem_mem_addr[5]), .A3(n141), .A4(
        ex_mem_addr[5]), .Y(n87) );
  AO22X1_LVT U41 ( .A1(n137), .A2(mem_mem_addr[4]), .A3(n141), .A4(
        ex_mem_addr[4]), .Y(n86) );
  AO22X1_LVT U42 ( .A1(n137), .A2(mem_mem_addr[3]), .A3(n141), .A4(
        ex_mem_addr[3]), .Y(n85) );
  AO22X1_LVT U43 ( .A1(n137), .A2(mem_mem_addr[2]), .A3(n141), .A4(
        ex_mem_addr[2]), .Y(n84) );
  AO22X1_LVT U48 ( .A1(n138), .A2(mem_mem_addr[1]), .A3(n141), .A4(
        ex_mem_addr[1]), .Y(n83) );
  AO22X1_LVT U49 ( .A1(n139), .A2(mem_mem_addr[0]), .A3(n143), .A4(
        ex_mem_addr[0]), .Y(n82) );
  AO22X1_LVT U50 ( .A1(n139), .A2(mem_aluop[4]), .A3(n143), .A4(ex_aluop[4]), 
        .Y(n78) );
  AO22X1_LVT U51 ( .A1(n138), .A2(mem_aluop[3]), .A3(n141), .A4(ex_aluop[3]), 
        .Y(n77) );
  AO22X1_LVT U52 ( .A1(n139), .A2(mem_aluop[2]), .A3(n143), .A4(ex_aluop[2]), 
        .Y(n76) );
  AO22X1_LVT U53 ( .A1(n138), .A2(mem_aluop[1]), .A3(n141), .A4(ex_aluop[1]), 
        .Y(n75) );
  AO22X1_LVT U54 ( .A1(n138), .A2(mem_aluop[0]), .A3(n141), .A4(ex_aluop[0]), 
        .Y(n74) );
  AO22X1_LVT U55 ( .A1(n138), .A2(mem_rt_data[31]), .A3(n141), .A4(
        ex_rt_data[31]), .Y(n73) );
  AO22X1_LVT U56 ( .A1(n138), .A2(mem_rt_data[30]), .A3(n141), .A4(
        ex_rt_data[30]), .Y(n72) );
  AO22X1_LVT U57 ( .A1(n138), .A2(mem_rt_data[29]), .A3(n141), .A4(
        ex_rt_data[29]), .Y(n71) );
  AO22X1_LVT U58 ( .A1(n139), .A2(mem_rt_data[28]), .A3(n143), .A4(
        ex_rt_data[28]), .Y(n70) );
  AO22X1_LVT U59 ( .A1(n139), .A2(mem_rt_data[27]), .A3(n143), .A4(
        ex_rt_data[27]), .Y(n69) );
  AO22X1_LVT U60 ( .A1(n139), .A2(mem_rt_data[26]), .A3(n143), .A4(
        ex_rt_data[26]), .Y(n68) );
  AO22X1_LVT U61 ( .A1(n139), .A2(mem_rt_data[25]), .A3(n143), .A4(
        ex_rt_data[25]), .Y(n67) );
  AO22X1_LVT U62 ( .A1(n139), .A2(mem_rt_data[24]), .A3(n143), .A4(
        ex_rt_data[24]), .Y(n66) );
  AO22X1_LVT U65 ( .A1(n139), .A2(mem_rt_data[23]), .A3(n143), .A4(
        ex_rt_data[23]), .Y(n65) );
  AO22X1_LVT U66 ( .A1(n139), .A2(mem_rt_data[22]), .A3(n143), .A4(
        ex_rt_data[22]), .Y(n64) );
  AO22X1_LVT U67 ( .A1(n139), .A2(mem_rt_data[21]), .A3(n143), .A4(
        ex_rt_data[21]), .Y(n63) );
  AO22X1_LVT U68 ( .A1(n139), .A2(mem_rt_data[20]), .A3(n143), .A4(
        ex_rt_data[20]), .Y(n62) );
  AO22X1_LVT U69 ( .A1(n139), .A2(mem_rt_data[19]), .A3(n143), .A4(
        ex_rt_data[19]), .Y(n61) );
  AO22X1_LVT U70 ( .A1(n139), .A2(mem_rt_data[18]), .A3(n143), .A4(
        ex_rt_data[18]), .Y(n60) );
  AO22X1_LVT U71 ( .A1(n139), .A2(mem_rt_data[17]), .A3(n143), .A4(
        ex_rt_data[17]), .Y(n59) );
  AO22X1_LVT U72 ( .A1(n139), .A2(mem_rt_data[16]), .A3(n143), .A4(
        ex_rt_data[16]), .Y(n58) );
  AO22X1_LVT U73 ( .A1(n139), .A2(mem_rt_data[15]), .A3(n143), .A4(
        ex_rt_data[15]), .Y(n57) );
  AO22X1_LVT U74 ( .A1(n139), .A2(mem_rt_data[14]), .A3(n143), .A4(
        ex_rt_data[14]), .Y(n56) );
  AO22X1_LVT U75 ( .A1(n139), .A2(mem_rt_data[13]), .A3(n143), .A4(
        ex_rt_data[13]), .Y(n55) );
  AO22X1_LVT U76 ( .A1(n139), .A2(mem_rt_data[12]), .A3(n143), .A4(
        ex_rt_data[12]), .Y(n54) );
  AO22X1_LVT U77 ( .A1(n139), .A2(mem_rt_data[11]), .A3(n143), .A4(
        ex_rt_data[11]), .Y(n53) );
  AO22X1_LVT U78 ( .A1(n139), .A2(mem_rt_data[10]), .A3(n143), .A4(
        ex_rt_data[10]), .Y(n52) );
  AO22X1_LVT U79 ( .A1(n139), .A2(mem_rt_data[9]), .A3(n143), .A4(
        ex_rt_data[9]), .Y(n51) );
  AO22X1_LVT U82 ( .A1(n139), .A2(mem_rt_data[8]), .A3(n143), .A4(
        ex_rt_data[8]), .Y(n50) );
  AO22X1_LVT U83 ( .A1(n139), .A2(mem_rt_data[7]), .A3(n143), .A4(
        ex_rt_data[7]), .Y(n49) );
  AO22X1_LVT U84 ( .A1(n139), .A2(mem_rt_data[6]), .A3(n143), .A4(
        ex_rt_data[6]), .Y(n48) );
  AO22X1_LVT U85 ( .A1(n139), .A2(mem_rt_data[5]), .A3(n143), .A4(
        ex_rt_data[5]), .Y(n47) );
  AO22X1_LVT U86 ( .A1(n138), .A2(mem_rt_data[4]), .A3(n141), .A4(
        ex_rt_data[4]), .Y(n46) );
  AO22X1_LVT U87 ( .A1(n138), .A2(mem_rt_data[3]), .A3(n141), .A4(
        ex_rt_data[3]), .Y(n45) );
  AO22X1_LVT U88 ( .A1(n138), .A2(mem_rt_data[2]), .A3(n141), .A4(
        ex_rt_data[2]), .Y(n44) );
  AO22X1_LVT U89 ( .A1(n138), .A2(mem_rt_data[1]), .A3(n141), .A4(
        ex_rt_data[1]), .Y(n43) );
  AO22X1_LVT U90 ( .A1(n138), .A2(mem_rt_data[0]), .A3(n141), .A4(
        ex_rt_data[0]), .Y(n42) );
  AO22X1_LVT U91 ( .A1(n138), .A2(mem_reg_waddr[4]), .A3(n141), .A4(
        ex_reg_waddr[4]), .Y(n41) );
  AO22X1_LVT U92 ( .A1(n138), .A2(mem_reg_waddr[3]), .A3(n141), .A4(
        ex_reg_waddr[3]), .Y(n40) );
  AO22X1_LVT U93 ( .A1(n138), .A2(mem_reg_waddr[2]), .A3(n141), .A4(
        ex_reg_waddr[2]), .Y(n39) );
  AO22X1_LVT U94 ( .A1(n138), .A2(mem_reg_waddr[1]), .A3(n141), .A4(
        ex_reg_waddr[1]), .Y(n38) );
  AO22X1_LVT U95 ( .A1(n138), .A2(mem_reg_waddr[0]), .A3(n141), .A4(
        ex_reg_waddr[0]), .Y(n37) );
  AO22X1_LVT U96 ( .A1(n138), .A2(mem_we), .A3(n141), .A4(ex_we), .Y(n36) );
  AO22X1_LVT U101 ( .A1(n136), .A2(mem_reg_wdata[31]), .A3(n140), .A4(
        ex_reg_wdata[31]), .Y(n35) );
  AO22X1_LVT U102 ( .A1(n136), .A2(mem_reg_wdata[30]), .A3(n140), .A4(
        ex_reg_wdata[30]), .Y(n34) );
  AO22X1_LVT U103 ( .A1(n136), .A2(mem_reg_wdata[29]), .A3(n140), .A4(
        ex_reg_wdata[29]), .Y(n33) );
  AO22X1_LVT U104 ( .A1(n136), .A2(mem_reg_wdata[28]), .A3(n140), .A4(
        ex_reg_wdata[28]), .Y(n32) );
  AO22X1_LVT U105 ( .A1(n136), .A2(mem_reg_wdata[27]), .A3(n140), .A4(
        ex_reg_wdata[27]), .Y(n31) );
  AO22X1_LVT U106 ( .A1(n136), .A2(mem_reg_wdata[26]), .A3(n140), .A4(
        ex_reg_wdata[26]), .Y(n30) );
  AO22X1_LVT U107 ( .A1(n136), .A2(mem_reg_wdata[25]), .A3(n140), .A4(
        ex_reg_wdata[25]), .Y(n29) );
  AO22X1_LVT U108 ( .A1(n136), .A2(mem_reg_wdata[24]), .A3(n140), .A4(
        ex_reg_wdata[24]), .Y(n28) );
  AO22X1_LVT U109 ( .A1(n136), .A2(mem_reg_wdata[23]), .A3(n140), .A4(
        ex_reg_wdata[23]), .Y(n27) );
  AO22X1_LVT U110 ( .A1(n136), .A2(mem_reg_wdata[22]), .A3(n140), .A4(
        ex_reg_wdata[22]), .Y(n26) );
  AO22X1_LVT U111 ( .A1(n136), .A2(mem_reg_wdata[21]), .A3(n140), .A4(
        ex_reg_wdata[21]), .Y(n25) );
  AO22X1_LVT U112 ( .A1(n136), .A2(mem_reg_wdata[20]), .A3(n140), .A4(
        ex_reg_wdata[20]), .Y(n24) );
  AO22X1_LVT U113 ( .A1(n136), .A2(mem_reg_wdata[19]), .A3(n140), .A4(
        ex_reg_wdata[19]), .Y(n23) );
  AO22X1_LVT U114 ( .A1(n136), .A2(mem_reg_wdata[18]), .A3(n140), .A4(
        ex_reg_wdata[18]), .Y(n22) );
  AO22X1_LVT U115 ( .A1(n136), .A2(mem_reg_wdata[17]), .A3(n140), .A4(
        ex_reg_wdata[17]), .Y(n21) );
  AO22X1_LVT U118 ( .A1(n136), .A2(mem_reg_wdata[16]), .A3(n140), .A4(
        ex_reg_wdata[16]), .Y(n20) );
  AO22X1_LVT U119 ( .A1(n136), .A2(mem_reg_wdata[15]), .A3(n140), .A4(
        ex_reg_wdata[15]), .Y(n19) );
  AO22X1_LVT U120 ( .A1(n136), .A2(mem_reg_wdata[14]), .A3(n140), .A4(
        ex_reg_wdata[14]), .Y(n18) );
  AO22X1_LVT U121 ( .A1(n136), .A2(mem_reg_wdata[13]), .A3(n140), .A4(
        ex_reg_wdata[13]), .Y(n17) );
  AO22X1_LVT U122 ( .A1(n136), .A2(mem_reg_wdata[12]), .A3(n140), .A4(
        ex_reg_wdata[12]), .Y(n16) );
  AO22X1_LVT U123 ( .A1(n136), .A2(mem_reg_wdata[11]), .A3(n140), .A4(
        ex_reg_wdata[11]), .Y(n15) );
  AO22X1_LVT U124 ( .A1(n136), .A2(mem_reg_wdata[10]), .A3(n140), .A4(
        ex_reg_wdata[10]), .Y(n14) );
  AO22X1_LVT U125 ( .A1(n136), .A2(mem_reg_wdata[9]), .A3(n140), .A4(
        ex_reg_wdata[9]), .Y(n13) );
  AO22X1_LVT U126 ( .A1(n136), .A2(mem_reg_wdata[8]), .A3(n140), .A4(
        ex_reg_wdata[8]), .Y(n12) );
  AO22X1_LVT U127 ( .A1(n136), .A2(mem_reg_wdata[7]), .A3(n140), .A4(
        ex_reg_wdata[7]), .Y(n11) );
  AO22X1_LVT U128 ( .A1(n136), .A2(mem_reg_wdata[6]), .A3(n140), .A4(
        ex_reg_wdata[6]), .Y(n10) );
  AO22X1_LVT U129 ( .A1(n136), .A2(mem_reg_wdata[5]), .A3(n140), .A4(
        ex_reg_wdata[5]), .Y(n9) );
  AO22X1_LVT U130 ( .A1(n136), .A2(mem_reg_wdata[4]), .A3(n140), .A4(
        ex_reg_wdata[4]), .Y(n8) );
  AO22X1_LVT U131 ( .A1(n136), .A2(mem_reg_wdata[3]), .A3(n140), .A4(
        ex_reg_wdata[3]), .Y(n7) );
  AO22X1_LVT U132 ( .A1(n136), .A2(mem_reg_wdata[2]), .A3(n140), .A4(
        ex_reg_wdata[2]), .Y(n6) );
  AO22X1_LVT U135 ( .A1(n136), .A2(mem_reg_wdata[1]), .A3(n140), .A4(
        ex_reg_wdata[1]), .Y(n5) );
  AO22X1_LVT U136 ( .A1(n136), .A2(mem_reg_wdata[0]), .A3(n140), .A4(
        ex_reg_wdata[0]), .Y(n4) );
  NOR2X0_LVT U8 ( .A1(stall[3]), .A2(rst), .Y(n3) );
  AND3X1_LVT U4 ( .A1(stall[3]), .A2(stall[4]), .A3(n135), .Y(n2) );
  INVX1_LVT U3 ( .A(rst), .Y(n135) );
  NBUFFX4_LVT U5 ( .A(n2), .Y(n136) );
  NBUFFX8_LVT U6 ( .A(n138), .Y(n137) );
  NBUFFX4_LVT U7 ( .A(n2), .Y(n138) );
  NBUFFX4_LVT U9 ( .A(n2), .Y(n139) );
  NBUFFX4_LVT U10 ( .A(n3), .Y(n140) );
  NBUFFX8_LVT U11 ( .A(n3), .Y(n141) );
  NBUFFX4_LVT U28 ( .A(n3), .Y(n143) );
  DFFX2_LVT \mem_aluop_reg[0]  ( .D(n74), .CLK(clk), .Q(mem_aluop[0]) );
  DFFX2_LVT \mem_aluop_reg[1]  ( .D(n75), .CLK(clk), .Q(mem_aluop[1]) );
  DFFX2_LVT \mem_mem_addr_reg[1]  ( .D(n83), .CLK(clk), .Q(mem_mem_addr[1]) );
  DFFX2_LVT \mem_rt_data_reg[2]  ( .D(n44), .CLK(clk), .Q(mem_rt_data[2]) );
  DFFX2_LVT \mem_rt_data_reg[3]  ( .D(n45), .CLK(clk), .Q(mem_rt_data[3]) );
  DFFX2_LVT \mem_rt_data_reg[1]  ( .D(n43), .CLK(clk), .Q(mem_rt_data[1]) );
  DFFX2_LVT \mem_rt_data_reg[4]  ( .D(n46), .CLK(clk), .Q(mem_rt_data[4]) );
endmodule


module stage_mem ( rst, reg_waddr_i, we_i, reg_wdata_i, mem_addr_i, aluop, 
        rt_data, mem_data_i, mem_busy, mem_done, reg_waddr_o, we_o, 
        reg_wdata_o, mem_addr_o, mem_re, mem_we, mem_sel, mem_data_o, stallreq
 );
  input [4:0] reg_waddr_i;
  input [31:0] reg_wdata_i;
  input [31:0] mem_addr_i;
  input [7:0] aluop;
  input [31:0] rt_data;
  input [31:0] mem_data_i;
  input [1:0] mem_busy;
  input [1:0] mem_done;
  output [4:0] reg_waddr_o;
  output [31:0] reg_wdata_o;
  output [31:0] mem_addr_o;
  output [3:0] mem_sel;
  output [31:0] mem_data_o;
  input rst, we_i;
  output we_o, mem_re, mem_we, stallreq;
  wire   mem_taking, N419, N420, N421, N422, N423, N424, N425, N426, N427,
         N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438,
         N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471,
         N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482,
         N483, N484, N485, N486, N487, N488, N489, N490, N492, N493, N494,
         N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505,
         N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516,
         N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527,
         N528, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n61, n63, n64, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n142, n143, n144, n145, n147, n150, n151, n152,
         n153, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n166, n167, n168, n170, n172, n174, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196;

  LATCHX1_LVT mem_taking_reg ( .CLK(N528), .D(N419), .Q(mem_taking) );
  LATCHX1_LVT we_o_reg ( .CLK(n191), .D(N490), .Q(we_o) );
  LATCHX1_LVT \mem_sel_reg[0]  ( .CLK(n190), .D(N524), .Q(mem_sel[0]) );
  LATCHX1_LVT \mem_sel_reg[1]  ( .CLK(n190), .D(N525), .Q(mem_sel[1]) );
  LATCHX1_LVT \mem_sel_reg[2]  ( .CLK(n190), .D(N526), .Q(mem_sel[2]) );
  LATCHX1_LVT \mem_sel_reg[3]  ( .CLK(n190), .D(N527), .Q(mem_sel[3]) );
  LATCHX1_LVT \mem_addr_o_reg[1]  ( .CLK(n191), .D(N422), .Q(mem_addr_o[1]) );
  LATCHX1_LVT \mem_addr_o_reg[2]  ( .CLK(n191), .D(N423), .Q(mem_addr_o[2]) );
  LATCHX1_LVT \mem_addr_o_reg[3]  ( .CLK(n191), .D(N424), .Q(mem_addr_o[3]) );
  LATCHX1_LVT \mem_addr_o_reg[4]  ( .CLK(n191), .D(N425), .Q(mem_addr_o[4]) );
  LATCHX1_LVT \mem_addr_o_reg[5]  ( .CLK(n191), .D(N426), .Q(mem_addr_o[5]) );
  LATCHX1_LVT \mem_addr_o_reg[6]  ( .CLK(n191), .D(N427), .Q(mem_addr_o[6]) );
  LATCHX1_LVT \mem_addr_o_reg[7]  ( .CLK(n191), .D(N428), .Q(mem_addr_o[7]) );
  LATCHX1_LVT \mem_addr_o_reg[8]  ( .CLK(n191), .D(N429), .Q(mem_addr_o[8]) );
  LATCHX1_LVT \mem_addr_o_reg[9]  ( .CLK(n191), .D(N430), .Q(mem_addr_o[9]) );
  LATCHX1_LVT \mem_addr_o_reg[10]  ( .CLK(n191), .D(N431), .Q(mem_addr_o[10])
         );
  LATCHX1_LVT \mem_addr_o_reg[11]  ( .CLK(n191), .D(N432), .Q(mem_addr_o[11])
         );
  LATCHX1_LVT \mem_addr_o_reg[12]  ( .CLK(n191), .D(N433), .Q(mem_addr_o[12])
         );
  LATCHX1_LVT \mem_addr_o_reg[13]  ( .CLK(n191), .D(N434), .Q(mem_addr_o[13])
         );
  LATCHX1_LVT \mem_addr_o_reg[14]  ( .CLK(n191), .D(N435), .Q(mem_addr_o[14])
         );
  LATCHX1_LVT \mem_addr_o_reg[15]  ( .CLK(n191), .D(N436), .Q(mem_addr_o[15])
         );
  LATCHX1_LVT \mem_addr_o_reg[16]  ( .CLK(n191), .D(N437), .Q(mem_addr_o[16])
         );
  LATCHX1_LVT \mem_addr_o_reg[17]  ( .CLK(n191), .D(N438), .Q(mem_addr_o[17])
         );
  LATCHX1_LVT \mem_addr_o_reg[18]  ( .CLK(n191), .D(N439), .Q(mem_addr_o[18])
         );
  LATCHX1_LVT \mem_addr_o_reg[19]  ( .CLK(n191), .D(N440), .Q(mem_addr_o[19])
         );
  LATCHX1_LVT \mem_addr_o_reg[20]  ( .CLK(n191), .D(N441), .Q(mem_addr_o[20])
         );
  LATCHX1_LVT \mem_addr_o_reg[21]  ( .CLK(n191), .D(N442), .Q(mem_addr_o[21])
         );
  LATCHX1_LVT \mem_addr_o_reg[22]  ( .CLK(n191), .D(N443), .Q(mem_addr_o[22])
         );
  LATCHX1_LVT \mem_addr_o_reg[23]  ( .CLK(n191), .D(N444), .Q(mem_addr_o[23])
         );
  LATCHX1_LVT \mem_addr_o_reg[24]  ( .CLK(n191), .D(N445), .Q(mem_addr_o[24])
         );
  LATCHX1_LVT \mem_addr_o_reg[25]  ( .CLK(n191), .D(N446), .Q(mem_addr_o[25])
         );
  LATCHX1_LVT \mem_addr_o_reg[26]  ( .CLK(n191), .D(N447), .Q(mem_addr_o[26])
         );
  LATCHX1_LVT \mem_addr_o_reg[27]  ( .CLK(n191), .D(N448), .Q(mem_addr_o[27])
         );
  LATCHX1_LVT \mem_addr_o_reg[28]  ( .CLK(n191), .D(N449), .Q(mem_addr_o[28])
         );
  LATCHX1_LVT \mem_addr_o_reg[29]  ( .CLK(n191), .D(N450), .Q(mem_addr_o[29])
         );
  LATCHX1_LVT \mem_addr_o_reg[30]  ( .CLK(n191), .D(N451), .Q(mem_addr_o[30])
         );
  LATCHX1_LVT \mem_addr_o_reg[31]  ( .CLK(n191), .D(N452), .Q(mem_addr_o[31])
         );
  LATCHX1_LVT \reg_wdata_o_reg[0]  ( .CLK(n196), .D(N492), .Q(reg_wdata_o[0])
         );
  LATCHX1_LVT \reg_wdata_o_reg[31]  ( .CLK(n196), .D(N523), .Q(reg_wdata_o[31]) );
  LATCHX1_LVT \reg_wdata_o_reg[30]  ( .CLK(n196), .D(N522), .Q(reg_wdata_o[30]) );
  LATCHX1_LVT \reg_wdata_o_reg[29]  ( .CLK(n196), .D(N521), .Q(reg_wdata_o[29]) );
  LATCHX1_LVT \reg_wdata_o_reg[28]  ( .CLK(n196), .D(N520), .Q(reg_wdata_o[28]) );
  LATCHX1_LVT \reg_wdata_o_reg[27]  ( .CLK(n196), .D(N519), .Q(reg_wdata_o[27]) );
  LATCHX1_LVT \reg_wdata_o_reg[26]  ( .CLK(n196), .D(N518), .Q(reg_wdata_o[26]) );
  LATCHX1_LVT \reg_wdata_o_reg[25]  ( .CLK(n196), .D(N517), .Q(reg_wdata_o[25]) );
  LATCHX1_LVT \reg_wdata_o_reg[24]  ( .CLK(n196), .D(N516), .Q(reg_wdata_o[24]) );
  LATCHX1_LVT \reg_wdata_o_reg[23]  ( .CLK(n196), .D(N515), .Q(reg_wdata_o[23]) );
  LATCHX1_LVT \reg_wdata_o_reg[22]  ( .CLK(n196), .D(N514), .Q(reg_wdata_o[22]) );
  LATCHX1_LVT \reg_wdata_o_reg[21]  ( .CLK(n196), .D(N513), .Q(reg_wdata_o[21]) );
  LATCHX1_LVT \reg_wdata_o_reg[20]  ( .CLK(n196), .D(N512), .Q(reg_wdata_o[20]) );
  LATCHX1_LVT \reg_wdata_o_reg[19]  ( .CLK(n196), .D(N511), .Q(reg_wdata_o[19]) );
  LATCHX1_LVT \reg_wdata_o_reg[18]  ( .CLK(n196), .D(N510), .Q(reg_wdata_o[18]) );
  LATCHX1_LVT \reg_wdata_o_reg[17]  ( .CLK(n196), .D(N509), .Q(reg_wdata_o[17]) );
  LATCHX1_LVT \reg_wdata_o_reg[16]  ( .CLK(n196), .D(N508), .Q(reg_wdata_o[16]) );
  LATCHX1_LVT \reg_wdata_o_reg[15]  ( .CLK(n196), .D(N507), .Q(reg_wdata_o[15]) );
  LATCHX1_LVT \reg_wdata_o_reg[14]  ( .CLK(n196), .D(N506), .Q(reg_wdata_o[14]) );
  LATCHX1_LVT \reg_wdata_o_reg[13]  ( .CLK(n196), .D(N505), .Q(reg_wdata_o[13]) );
  LATCHX1_LVT \reg_wdata_o_reg[12]  ( .CLK(n196), .D(N504), .Q(reg_wdata_o[12]) );
  LATCHX1_LVT \reg_wdata_o_reg[11]  ( .CLK(n196), .D(N503), .Q(reg_wdata_o[11]) );
  LATCHX1_LVT \reg_wdata_o_reg[10]  ( .CLK(n11), .D(N502), .Q(reg_wdata_o[10])
         );
  LATCHX1_LVT \reg_wdata_o_reg[9]  ( .CLK(n11), .D(N501), .Q(reg_wdata_o[9])
         );
  LATCHX1_LVT \reg_wdata_o_reg[8]  ( .CLK(n196), .D(N500), .Q(reg_wdata_o[8])
         );
  LATCHX1_LVT \reg_wdata_o_reg[7]  ( .CLK(n196), .D(N499), .Q(reg_wdata_o[7])
         );
  LATCHX1_LVT \reg_wdata_o_reg[6]  ( .CLK(n196), .D(N498), .Q(reg_wdata_o[6])
         );
  LATCHX1_LVT \reg_wdata_o_reg[5]  ( .CLK(n11), .D(N497), .Q(reg_wdata_o[5])
         );
  LATCHX1_LVT \reg_wdata_o_reg[4]  ( .CLK(n11), .D(N496), .Q(reg_wdata_o[4])
         );
  LATCHX1_LVT \reg_wdata_o_reg[3]  ( .CLK(n196), .D(N495), .Q(reg_wdata_o[3])
         );
  LATCHX1_LVT \reg_wdata_o_reg[2]  ( .CLK(n196), .D(N494), .Q(reg_wdata_o[2])
         );
  LATCHX1_LVT \reg_wdata_o_reg[1]  ( .CLK(n196), .D(N493), .Q(reg_wdata_o[1])
         );
  LATCHX1_LVT mem_re_reg ( .CLK(n190), .D(N419), .Q(mem_re) );
  LATCHX1_LVT \reg_waddr_o_reg[4]  ( .CLK(n191), .D(N489), .Q(reg_waddr_o[4])
         );
  LATCHX1_LVT \reg_waddr_o_reg[3]  ( .CLK(n191), .D(N488), .Q(reg_waddr_o[3])
         );
  LATCHX1_LVT \reg_waddr_o_reg[2]  ( .CLK(n191), .D(N487), .Q(reg_waddr_o[2])
         );
  LATCHX1_LVT \reg_waddr_o_reg[1]  ( .CLK(n191), .D(N486), .Q(reg_waddr_o[1])
         );
  LATCHX1_LVT \reg_waddr_o_reg[0]  ( .CLK(n191), .D(N485), .Q(reg_waddr_o[0])
         );
  LATCHX1_LVT mem_we_reg ( .CLK(n190), .D(N420), .Q(mem_we) );
  LATCHX1_LVT \mem_data_o_reg[31]  ( .CLK(n190), .D(N484), .Q(mem_data_o[31])
         );
  LATCHX1_LVT \mem_data_o_reg[30]  ( .CLK(n190), .D(N483), .Q(mem_data_o[30])
         );
  LATCHX1_LVT \mem_data_o_reg[29]  ( .CLK(n190), .D(N482), .Q(mem_data_o[29])
         );
  LATCHX1_LVT \mem_data_o_reg[28]  ( .CLK(n190), .D(N481), .Q(mem_data_o[28])
         );
  LATCHX1_LVT \mem_data_o_reg[27]  ( .CLK(n190), .D(N480), .Q(mem_data_o[27])
         );
  LATCHX1_LVT \mem_data_o_reg[26]  ( .CLK(n190), .D(N479), .Q(mem_data_o[26])
         );
  LATCHX1_LVT \mem_data_o_reg[25]  ( .CLK(n190), .D(N478), .Q(mem_data_o[25])
         );
  LATCHX1_LVT \mem_data_o_reg[24]  ( .CLK(n190), .D(N477), .Q(mem_data_o[24])
         );
  LATCHX1_LVT \mem_data_o_reg[23]  ( .CLK(n190), .D(N476), .Q(mem_data_o[23])
         );
  LATCHX1_LVT \mem_data_o_reg[22]  ( .CLK(n190), .D(N475), .Q(mem_data_o[22])
         );
  LATCHX1_LVT \mem_data_o_reg[21]  ( .CLK(n190), .D(N474), .Q(mem_data_o[21])
         );
  LATCHX1_LVT \mem_data_o_reg[20]  ( .CLK(n190), .D(N473), .Q(mem_data_o[20])
         );
  LATCHX1_LVT \mem_data_o_reg[19]  ( .CLK(n190), .D(N472), .Q(mem_data_o[19])
         );
  LATCHX1_LVT \mem_data_o_reg[18]  ( .CLK(n190), .D(N471), .Q(mem_data_o[18])
         );
  LATCHX1_LVT \mem_data_o_reg[17]  ( .CLK(n190), .D(N470), .Q(mem_data_o[17])
         );
  LATCHX1_LVT \mem_data_o_reg[16]  ( .CLK(n190), .D(N469), .Q(mem_data_o[16])
         );
  LATCHX1_LVT \mem_data_o_reg[15]  ( .CLK(n190), .D(N468), .Q(mem_data_o[15])
         );
  LATCHX1_LVT \mem_data_o_reg[14]  ( .CLK(n190), .D(N467), .Q(mem_data_o[14])
         );
  LATCHX1_LVT \mem_data_o_reg[13]  ( .CLK(n190), .D(N466), .Q(mem_data_o[13])
         );
  LATCHX1_LVT \mem_data_o_reg[12]  ( .CLK(n190), .D(N465), .Q(mem_data_o[12])
         );
  LATCHX1_LVT \mem_data_o_reg[11]  ( .CLK(n190), .D(N464), .Q(mem_data_o[11])
         );
  LATCHX1_LVT \mem_data_o_reg[10]  ( .CLK(n190), .D(N463), .Q(mem_data_o[10])
         );
  LATCHX1_LVT \mem_data_o_reg[9]  ( .CLK(n190), .D(N462), .Q(mem_data_o[9]) );
  LATCHX1_LVT \mem_data_o_reg[8]  ( .CLK(n190), .D(N461), .Q(mem_data_o[8]) );
  LATCHX1_LVT \mem_data_o_reg[7]  ( .CLK(n190), .D(N460), .Q(mem_data_o[7]) );
  LATCHX1_LVT \mem_data_o_reg[6]  ( .CLK(n190), .D(N459), .Q(mem_data_o[6]) );
  LATCHX1_LVT \mem_data_o_reg[5]  ( .CLK(n190), .D(N458), .Q(mem_data_o[5]) );
  LATCHX1_LVT \mem_data_o_reg[4]  ( .CLK(n190), .D(N457), .Q(mem_data_o[4]) );
  LATCHX1_LVT \mem_data_o_reg[3]  ( .CLK(n190), .D(N456), .Q(mem_data_o[3]) );
  LATCHX1_LVT \mem_data_o_reg[2]  ( .CLK(n190), .D(N455), .Q(mem_data_o[2]) );
  LATCHX1_LVT \mem_data_o_reg[1]  ( .CLK(n190), .D(N454), .Q(mem_data_o[1]) );
  LATCHX1_LVT \mem_data_o_reg[0]  ( .CLK(n190), .D(N453), .Q(mem_data_o[0]) );
  OR2X1_LVT U3 ( .A1(mem_busy[1]), .A2(mem_busy[0]), .Y(n172) );
  OR3X2_LVT U4 ( .A1(rst), .A2(mem_taking), .A3(n172), .Y(n20) );
  AND2X1_LVT U6 ( .A1(aluop[4]), .A2(n189), .Y(n2) );
  INVX1_LVT U7 ( .A(aluop[3]), .Y(n1) );
  NAND2X0_LVT U8 ( .A1(aluop[2]), .A2(n1), .Y(n6) );
  OR2X1_LVT U11 ( .A1(n1), .A2(aluop[2]), .Y(n8) );
  INVX1_LVT U12 ( .A(n8), .Y(n7) );
  NAND3X0_LVT U13 ( .A1(n186), .A2(n185), .A3(n7), .Y(n16) );
  NAND2X0_LVT U14 ( .A1(n6), .A2(n16), .Y(n17) );
  NAND2X0_LVT U15 ( .A1(n2), .A2(n17), .Y(n174) );
  INVX1_LVT U16 ( .A(n174), .Y(N419) );
  NAND4X0_LVT U17 ( .A1(aluop[4]), .A2(n7), .A3(n189), .A4(aluop[1]), .Y(n145)
         );
  NAND4X0_LVT U18 ( .A1(n7), .A2(aluop[0]), .A3(n2), .A4(n186), .Y(n150) );
  OR3X1_LVT U21 ( .A1(mem_taking), .A2(mem_busy[1]), .A3(mem_busy[0]), .Y(n3)
         );
  NAND2X0_LVT U22 ( .A1(n184), .A2(n3), .Y(n4) );
  INVX1_LVT U27 ( .A(n172), .Y(n5) );
  NAND2X0_LVT U28 ( .A1(mem_taking), .A2(n5), .Y(n15) );
  INVX1_LVT U29 ( .A(n6), .Y(n59) );
  OA21X1_LVT U30 ( .A1(n7), .A2(n59), .A3(aluop[4]), .Y(n21) );
  AND2X1_LVT U31 ( .A1(n186), .A2(n185), .Y(n9) );
  AO221X1_LVT U32 ( .A1(n21), .A2(n9), .A3(n21), .A4(n8), .A5(n20), .Y(n10) );
  INVX1_LVT U42 ( .A(n15), .Y(n18) );
  NAND3X0_LVT U43 ( .A1(aluop[4]), .A2(n18), .A3(n184), .Y(n120) );
  INVX2_LVT U44 ( .A(n120), .Y(n119) );
  AND2X1_LVT U47 ( .A1(n188), .A2(n187), .Y(n151) );
  NAND3X0_LVT U48 ( .A1(n59), .A2(aluop[0]), .A3(n186), .Y(n121) );
  NAND2X0_LVT U49 ( .A1(n16), .A2(n121), .Y(n70) );
  AND4X1_LVT U50 ( .A1(aluop[1]), .A2(n59), .A3(n151), .A4(n185), .Y(n118) );
  AO21X1_LVT U51 ( .A1(n151), .A2(n70), .A3(n118), .Y(n67) );
  AND2X1_LVT U52 ( .A1(n119), .A2(n67), .Y(n57) );
  INVX1_LVT U53 ( .A(n17), .Y(n109) );
  NAND2X0_LVT U54 ( .A1(n18), .A2(n184), .Y(n19) );
  OAI22X1_LVT U55 ( .A1(n21), .A2(n20), .A3(aluop[4]), .A4(n19), .Y(n116) );
  AO22X1_LVT U58 ( .A1(mem_data_i[15]), .A2(n57), .A3(reg_wdata_i[15]), .A4(
        n194), .Y(n22) );
  INVX1_LVT U59 ( .A(n22), .Y(n27) );
  OA221X1_LVT U60 ( .A1(mem_addr_i[1]), .A2(mem_data_i[15]), .A3(n188), .A4(
        mem_data_i[31]), .A5(mem_addr_i[0]), .Y(n24) );
  AND2X1_LVT U61 ( .A1(mem_addr_i[1]), .A2(n187), .Y(n147) );
  AO22X1_LVT U62 ( .A1(n147), .A2(mem_data_i[23]), .A3(n151), .A4(
        mem_data_i[7]), .Y(n23) );
  OR2X1_LVT U63 ( .A1(n24), .A2(n23), .Y(n61) );
  NAND4X0_LVT U64 ( .A1(n59), .A2(n185), .A3(n186), .A4(n61), .Y(n123) );
  NOR2X2_LVT U65 ( .A1(n120), .A2(n123), .Y(n53) );
  INVX1_LVT U66 ( .A(n53), .Y(n26) );
  AND3X1_LVT U67 ( .A1(n147), .A2(n119), .A3(n70), .Y(n63) );
  NAND2X0_LVT U68 ( .A1(n63), .A2(mem_data_i[31]), .Y(n25) );
  NAND3X0_LVT U69 ( .A1(n27), .A2(n26), .A3(n25), .Y(N507) );
  AO22X1_LVT U70 ( .A1(mem_data_i[30]), .A2(n63), .A3(reg_wdata_i[14]), .A4(
        n194), .Y(n28) );
  INVX1_LVT U71 ( .A(n28), .Y(n31) );
  INVX1_LVT U72 ( .A(n53), .Y(n30) );
  NAND2X0_LVT U73 ( .A1(n57), .A2(mem_data_i[14]), .Y(n29) );
  NAND3X0_LVT U74 ( .A1(n31), .A2(n30), .A3(n29), .Y(N506) );
  AO22X1_LVT U75 ( .A1(mem_data_i[29]), .A2(n63), .A3(reg_wdata_i[13]), .A4(
        n194), .Y(n32) );
  INVX1_LVT U76 ( .A(n32), .Y(n35) );
  INVX1_LVT U77 ( .A(n53), .Y(n34) );
  NAND2X0_LVT U78 ( .A1(n57), .A2(mem_data_i[13]), .Y(n33) );
  NAND3X0_LVT U79 ( .A1(n35), .A2(n34), .A3(n33), .Y(N505) );
  AO22X1_LVT U80 ( .A1(mem_data_i[28]), .A2(n63), .A3(reg_wdata_i[12]), .A4(
        n194), .Y(n36) );
  INVX1_LVT U81 ( .A(n36), .Y(n39) );
  INVX1_LVT U82 ( .A(n53), .Y(n38) );
  NAND2X0_LVT U83 ( .A1(n57), .A2(mem_data_i[12]), .Y(n37) );
  NAND3X0_LVT U84 ( .A1(n39), .A2(n38), .A3(n37), .Y(N504) );
  AO22X1_LVT U85 ( .A1(mem_data_i[27]), .A2(n63), .A3(reg_wdata_i[11]), .A4(
        n194), .Y(n40) );
  INVX1_LVT U86 ( .A(n40), .Y(n43) );
  INVX1_LVT U87 ( .A(n53), .Y(n42) );
  NAND2X0_LVT U88 ( .A1(n57), .A2(mem_data_i[11]), .Y(n41) );
  NAND3X0_LVT U89 ( .A1(n43), .A2(n42), .A3(n41), .Y(N503) );
  AO22X1_LVT U90 ( .A1(mem_data_i[26]), .A2(n63), .A3(reg_wdata_i[10]), .A4(
        n194), .Y(n44) );
  INVX1_LVT U91 ( .A(n44), .Y(n47) );
  INVX1_LVT U92 ( .A(n53), .Y(n46) );
  NAND2X0_LVT U93 ( .A1(n57), .A2(mem_data_i[10]), .Y(n45) );
  NAND3X0_LVT U94 ( .A1(n47), .A2(n46), .A3(n45), .Y(N502) );
  AO22X1_LVT U95 ( .A1(mem_data_i[25]), .A2(n63), .A3(reg_wdata_i[9]), .A4(
        n194), .Y(n48) );
  INVX1_LVT U96 ( .A(n48), .Y(n51) );
  INVX1_LVT U97 ( .A(n53), .Y(n50) );
  NAND2X0_LVT U98 ( .A1(n57), .A2(mem_data_i[9]), .Y(n49) );
  NAND3X0_LVT U99 ( .A1(n51), .A2(n50), .A3(n49), .Y(N501) );
  AO22X1_LVT U100 ( .A1(mem_data_i[24]), .A2(n63), .A3(reg_wdata_i[8]), .A4(
        n194), .Y(n52) );
  INVX1_LVT U101 ( .A(n52), .Y(n56) );
  INVX1_LVT U102 ( .A(n53), .Y(n55) );
  NAND2X0_LVT U103 ( .A1(n57), .A2(mem_data_i[8]), .Y(n54) );
  NAND3X0_LVT U104 ( .A1(n56), .A2(n55), .A3(n54), .Y(N500) );
  AO22X1_LVT U105 ( .A1(mem_data_i[7]), .A2(n57), .A3(reg_wdata_i[7]), .A4(
        n194), .Y(n58) );
  INVX1_LVT U106 ( .A(n58), .Y(n66) );
  OA221X1_LVT U107 ( .A1(aluop[1]), .A2(n185), .A3(n186), .A4(aluop[0]), .A5(
        n59), .Y(n71) );
  NAND2X0_LVT U110 ( .A1(mem_data_i[23]), .A2(n63), .Y(n64) );
  NAND3X0_LVT U111 ( .A1(n66), .A2(n193), .A3(n64), .Y(N499) );
  AND3X1_LVT U112 ( .A1(mem_addr_i[0]), .A2(n71), .A3(n188), .Y(n107) );
  AO21X1_LVT U113 ( .A1(n71), .A2(n151), .A3(n67), .Y(n106) );
  AO22X1_LVT U114 ( .A1(mem_data_i[8]), .A2(n107), .A3(mem_data_i[0]), .A4(
        n106), .Y(n68) );
  INVX1_LVT U115 ( .A(n68), .Y(n74) );
  AND3X1_LVT U116 ( .A1(mem_addr_i[1]), .A2(mem_addr_i[0]), .A3(n71), .Y(n110)
         );
  AO22X1_LVT U117 ( .A1(reg_wdata_i[0]), .A2(n109), .A3(mem_data_i[24]), .A4(
        n110), .Y(n69) );
  INVX1_LVT U118 ( .A(n69), .Y(n73) );
  OA21X1_LVT U119 ( .A1(n71), .A2(n70), .A3(n147), .Y(n112) );
  NAND2X0_LVT U120 ( .A1(mem_data_i[16]), .A2(n112), .Y(n72) );
  NAND3X0_LVT U121 ( .A1(n74), .A2(n73), .A3(n72), .Y(n75) );
  AO22X1_LVT U122 ( .A1(n119), .A2(n75), .A3(reg_wdata_i[0]), .A4(n116), .Y(
        N492) );
  AO22X1_LVT U123 ( .A1(n107), .A2(mem_data_i[9]), .A3(mem_data_i[1]), .A4(
        n106), .Y(n76) );
  INVX1_LVT U124 ( .A(n76), .Y(n80) );
  AO22X1_LVT U125 ( .A1(n110), .A2(mem_data_i[25]), .A3(n109), .A4(
        reg_wdata_i[1]), .Y(n77) );
  INVX1_LVT U126 ( .A(n77), .Y(n79) );
  NAND2X0_LVT U127 ( .A1(n112), .A2(mem_data_i[17]), .Y(n78) );
  NAND3X0_LVT U128 ( .A1(n80), .A2(n79), .A3(n78), .Y(n81) );
  AO22X1_LVT U129 ( .A1(n119), .A2(n81), .A3(reg_wdata_i[1]), .A4(n116), .Y(
        N493) );
  AO22X1_LVT U130 ( .A1(n107), .A2(mem_data_i[10]), .A3(mem_data_i[2]), .A4(
        n106), .Y(n82) );
  INVX1_LVT U131 ( .A(n82), .Y(n86) );
  AO22X1_LVT U132 ( .A1(n110), .A2(mem_data_i[26]), .A3(n109), .A4(
        reg_wdata_i[2]), .Y(n83) );
  INVX1_LVT U133 ( .A(n83), .Y(n85) );
  NAND2X0_LVT U134 ( .A1(n112), .A2(mem_data_i[18]), .Y(n84) );
  NAND3X0_LVT U135 ( .A1(n86), .A2(n85), .A3(n84), .Y(n87) );
  AO22X1_LVT U136 ( .A1(n119), .A2(n87), .A3(reg_wdata_i[2]), .A4(n116), .Y(
        N494) );
  AO22X1_LVT U137 ( .A1(n107), .A2(mem_data_i[11]), .A3(mem_data_i[3]), .A4(
        n106), .Y(n88) );
  INVX1_LVT U138 ( .A(n88), .Y(n92) );
  AO22X1_LVT U139 ( .A1(n110), .A2(mem_data_i[27]), .A3(n109), .A4(
        reg_wdata_i[3]), .Y(n89) );
  INVX1_LVT U140 ( .A(n89), .Y(n91) );
  NAND2X0_LVT U141 ( .A1(n112), .A2(mem_data_i[19]), .Y(n90) );
  NAND3X0_LVT U142 ( .A1(n92), .A2(n91), .A3(n90), .Y(n93) );
  AO22X1_LVT U143 ( .A1(n119), .A2(n93), .A3(reg_wdata_i[3]), .A4(n116), .Y(
        N495) );
  AO22X1_LVT U144 ( .A1(n107), .A2(mem_data_i[12]), .A3(mem_data_i[4]), .A4(
        n106), .Y(n94) );
  INVX1_LVT U145 ( .A(n94), .Y(n98) );
  AO22X1_LVT U146 ( .A1(n110), .A2(mem_data_i[28]), .A3(n109), .A4(
        reg_wdata_i[4]), .Y(n95) );
  INVX1_LVT U147 ( .A(n95), .Y(n97) );
  NAND2X0_LVT U148 ( .A1(n112), .A2(mem_data_i[20]), .Y(n96) );
  NAND3X0_LVT U149 ( .A1(n98), .A2(n97), .A3(n96), .Y(n99) );
  AO22X1_LVT U150 ( .A1(n119), .A2(n99), .A3(reg_wdata_i[4]), .A4(n116), .Y(
        N496) );
  AO22X1_LVT U151 ( .A1(n107), .A2(mem_data_i[13]), .A3(mem_data_i[5]), .A4(
        n106), .Y(n100) );
  INVX1_LVT U152 ( .A(n100), .Y(n104) );
  AO22X1_LVT U153 ( .A1(n110), .A2(mem_data_i[29]), .A3(n109), .A4(
        reg_wdata_i[5]), .Y(n101) );
  INVX1_LVT U154 ( .A(n101), .Y(n103) );
  NAND2X0_LVT U155 ( .A1(n112), .A2(mem_data_i[21]), .Y(n102) );
  NAND3X0_LVT U156 ( .A1(n104), .A2(n103), .A3(n102), .Y(n105) );
  AO22X1_LVT U157 ( .A1(n119), .A2(n105), .A3(reg_wdata_i[5]), .A4(n116), .Y(
        N497) );
  AO22X1_LVT U158 ( .A1(n107), .A2(mem_data_i[14]), .A3(mem_data_i[6]), .A4(
        n106), .Y(n108) );
  INVX1_LVT U159 ( .A(n108), .Y(n115) );
  AO22X1_LVT U160 ( .A1(n110), .A2(mem_data_i[30]), .A3(n109), .A4(
        reg_wdata_i[6]), .Y(n111) );
  INVX1_LVT U161 ( .A(n111), .Y(n114) );
  NAND2X0_LVT U162 ( .A1(n112), .A2(mem_data_i[22]), .Y(n113) );
  NAND3X0_LVT U163 ( .A1(n115), .A2(n114), .A3(n113), .Y(n117) );
  AO22X1_LVT U164 ( .A1(n119), .A2(n117), .A3(reg_wdata_i[6]), .A4(n116), .Y(
        N498) );
  AND2X2_LVT U165 ( .A1(n119), .A2(n118), .Y(n142) );
  AOI22X1_LVT U166 ( .A1(mem_data_i[16]), .A2(n142), .A3(reg_wdata_i[16]), 
        .A4(n131), .Y(n124) );
  NAND2X0_LVT U167 ( .A1(mem_data_i[15]), .A2(n187), .Y(n122) );
  AO221X2_LVT U168 ( .A1(n123), .A2(n122), .A3(n123), .A4(n121), .A5(n120), 
        .Y(n143) );
  NAND2X0_LVT U169 ( .A1(n124), .A2(n143), .Y(N508) );
  AOI22X1_LVT U170 ( .A1(mem_data_i[17]), .A2(n142), .A3(reg_wdata_i[17]), 
        .A4(n194), .Y(n125) );
  NAND2X0_LVT U171 ( .A1(n125), .A2(n143), .Y(N509) );
  AOI22X1_LVT U172 ( .A1(mem_data_i[18]), .A2(n142), .A3(reg_wdata_i[18]), 
        .A4(n131), .Y(n126) );
  NAND2X0_LVT U173 ( .A1(n126), .A2(n143), .Y(N510) );
  AOI22X1_LVT U174 ( .A1(mem_data_i[19]), .A2(n142), .A3(reg_wdata_i[19]), 
        .A4(n131), .Y(n127) );
  NAND2X0_LVT U175 ( .A1(n127), .A2(n143), .Y(N511) );
  AOI22X1_LVT U176 ( .A1(mem_data_i[20]), .A2(n142), .A3(reg_wdata_i[20]), 
        .A4(n131), .Y(n128) );
  NAND2X0_LVT U177 ( .A1(n128), .A2(n143), .Y(N512) );
  AOI22X1_LVT U178 ( .A1(mem_data_i[21]), .A2(n142), .A3(reg_wdata_i[21]), 
        .A4(n131), .Y(n130) );
  NAND2X0_LVT U179 ( .A1(n130), .A2(n143), .Y(N513) );
  AOI22X1_LVT U181 ( .A1(mem_data_i[22]), .A2(n142), .A3(reg_wdata_i[22]), 
        .A4(n131), .Y(n132) );
  NAND2X0_LVT U182 ( .A1(n132), .A2(n143), .Y(N514) );
  AOI22X1_LVT U183 ( .A1(mem_data_i[23]), .A2(n142), .A3(reg_wdata_i[23]), 
        .A4(n131), .Y(n133) );
  NAND2X0_LVT U184 ( .A1(n133), .A2(n143), .Y(N515) );
  AOI22X1_LVT U185 ( .A1(mem_data_i[24]), .A2(n142), .A3(reg_wdata_i[24]), 
        .A4(n194), .Y(n134) );
  NAND2X0_LVT U186 ( .A1(n134), .A2(n143), .Y(N516) );
  AOI22X1_LVT U187 ( .A1(mem_data_i[25]), .A2(n142), .A3(reg_wdata_i[25]), 
        .A4(n131), .Y(n135) );
  NAND2X0_LVT U188 ( .A1(n135), .A2(n143), .Y(N517) );
  AOI22X1_LVT U189 ( .A1(mem_data_i[26]), .A2(n142), .A3(reg_wdata_i[26]), 
        .A4(n194), .Y(n136) );
  NAND2X0_LVT U190 ( .A1(n136), .A2(n143), .Y(N518) );
  AOI22X1_LVT U191 ( .A1(mem_data_i[27]), .A2(n142), .A3(reg_wdata_i[27]), 
        .A4(n194), .Y(n137) );
  NAND2X0_LVT U192 ( .A1(n137), .A2(n143), .Y(N519) );
  AOI22X1_LVT U193 ( .A1(mem_data_i[28]), .A2(n142), .A3(reg_wdata_i[28]), 
        .A4(n194), .Y(n138) );
  NAND2X0_LVT U194 ( .A1(n138), .A2(n143), .Y(N520) );
  AOI22X1_LVT U195 ( .A1(mem_data_i[29]), .A2(n142), .A3(reg_wdata_i[29]), 
        .A4(n194), .Y(n139) );
  NAND2X0_LVT U196 ( .A1(n139), .A2(n143), .Y(N521) );
  AOI22X1_LVT U197 ( .A1(mem_data_i[30]), .A2(n142), .A3(reg_wdata_i[30]), 
        .A4(n194), .Y(n140) );
  NAND2X0_LVT U198 ( .A1(n140), .A2(n143), .Y(N522) );
  AOI22X1_LVT U199 ( .A1(mem_data_i[31]), .A2(n142), .A3(reg_wdata_i[31]), 
        .A4(n194), .Y(n144) );
  NAND2X0_LVT U200 ( .A1(n144), .A2(n143), .Y(N523) );
  AND2X1_LVT U201 ( .A1(n151), .A2(N420), .Y(N524) );
  INVX2_LVT U202 ( .A(n145), .Y(n155) );
  OA221X1_LVT U204 ( .A1(mem_addr_i[0]), .A2(n155), .A3(n187), .A4(n192), .A5(
        n188), .Y(N525) );
  NAND2X0_LVT U205 ( .A1(n155), .A2(n185), .Y(n157) );
  NAND2X0_LVT U206 ( .A1(n150), .A2(n157), .Y(n156) );
  AND2X2_LVT U207 ( .A1(aluop[0]), .A2(n155), .Y(n166) );
  AO22X1_LVT U208 ( .A1(n147), .A2(n156), .A3(n151), .A4(n166), .Y(N526) );
  AO221X1_LVT U209 ( .A1(mem_addr_i[0]), .A2(n150), .A3(n187), .A4(n157), .A5(
        n188), .Y(n153) );
  NAND2X0_LVT U210 ( .A1(n151), .A2(n166), .Y(n152) );
  NAND2X0_LVT U211 ( .A1(n153), .A2(n152), .Y(N527) );
  AND2X1_LVT U212 ( .A1(n189), .A2(we_i), .Y(N490) );
  AND2X1_LVT U213 ( .A1(n189), .A2(reg_waddr_i[0]), .Y(N485) );
  AND2X1_LVT U214 ( .A1(n189), .A2(reg_waddr_i[1]), .Y(N486) );
  AND2X1_LVT U215 ( .A1(n189), .A2(reg_waddr_i[2]), .Y(N487) );
  AND2X1_LVT U216 ( .A1(n189), .A2(reg_waddr_i[3]), .Y(N488) );
  AND2X1_LVT U217 ( .A1(n189), .A2(reg_waddr_i[4]), .Y(N489) );
  AND2X1_LVT U218 ( .A1(rt_data[0]), .A2(N420), .Y(N453) );
  AND2X1_LVT U219 ( .A1(rt_data[1]), .A2(N420), .Y(N454) );
  AND2X1_LVT U220 ( .A1(rt_data[2]), .A2(N420), .Y(N455) );
  AND2X1_LVT U221 ( .A1(rt_data[3]), .A2(N420), .Y(N456) );
  AND2X1_LVT U222 ( .A1(rt_data[4]), .A2(N420), .Y(N457) );
  AND2X1_LVT U223 ( .A1(rt_data[5]), .A2(N420), .Y(N458) );
  AND2X1_LVT U224 ( .A1(rt_data[6]), .A2(N420), .Y(N459) );
  AND2X1_LVT U225 ( .A1(rt_data[7]), .A2(N420), .Y(N460) );
  AO22X1_LVT U226 ( .A1(n155), .A2(rt_data[8]), .A3(n192), .A4(rt_data[0]), 
        .Y(N461) );
  AO22X1_LVT U227 ( .A1(n155), .A2(rt_data[9]), .A3(n192), .A4(rt_data[1]), 
        .Y(N462) );
  AO22X1_LVT U228 ( .A1(n155), .A2(rt_data[10]), .A3(n192), .A4(rt_data[2]), 
        .Y(N463) );
  AO22X1_LVT U229 ( .A1(n155), .A2(rt_data[11]), .A3(n192), .A4(rt_data[3]), 
        .Y(N464) );
  AO22X1_LVT U230 ( .A1(n155), .A2(rt_data[12]), .A3(n192), .A4(rt_data[4]), 
        .Y(N465) );
  AO22X1_LVT U231 ( .A1(n155), .A2(rt_data[13]), .A3(n192), .A4(rt_data[5]), 
        .Y(N466) );
  AO22X1_LVT U232 ( .A1(n155), .A2(rt_data[14]), .A3(n192), .A4(rt_data[6]), 
        .Y(N467) );
  AO22X1_LVT U233 ( .A1(n155), .A2(rt_data[15]), .A3(n192), .A4(rt_data[7]), 
        .Y(N468) );
  AO22X1_LVT U234 ( .A1(n166), .A2(rt_data[16]), .A3(rt_data[0]), .A4(n156), 
        .Y(N469) );
  AO22X1_LVT U235 ( .A1(n166), .A2(rt_data[17]), .A3(rt_data[1]), .A4(n156), 
        .Y(N470) );
  AO22X1_LVT U236 ( .A1(n166), .A2(rt_data[18]), .A3(rt_data[2]), .A4(n156), 
        .Y(N471) );
  AO22X1_LVT U237 ( .A1(n166), .A2(rt_data[19]), .A3(rt_data[3]), .A4(n156), 
        .Y(N472) );
  AO22X1_LVT U238 ( .A1(n166), .A2(rt_data[20]), .A3(rt_data[4]), .A4(n156), 
        .Y(N473) );
  AO22X1_LVT U239 ( .A1(n166), .A2(rt_data[21]), .A3(rt_data[5]), .A4(n156), 
        .Y(N474) );
  AO22X1_LVT U240 ( .A1(n166), .A2(rt_data[22]), .A3(rt_data[6]), .A4(n156), 
        .Y(N475) );
  AO22X1_LVT U241 ( .A1(n166), .A2(rt_data[23]), .A3(rt_data[7]), .A4(n156), 
        .Y(N476) );
  INVX1_LVT U242 ( .A(n157), .Y(n168) );
  AO22X1_LVT U243 ( .A1(n166), .A2(rt_data[24]), .A3(n192), .A4(rt_data[0]), 
        .Y(n158) );
  AO21X1_LVT U244 ( .A1(n168), .A2(rt_data[8]), .A3(n158), .Y(N477) );
  AO22X1_LVT U245 ( .A1(n166), .A2(rt_data[25]), .A3(n192), .A4(rt_data[1]), 
        .Y(n159) );
  AO21X1_LVT U246 ( .A1(n168), .A2(rt_data[9]), .A3(n159), .Y(N478) );
  AO22X1_LVT U247 ( .A1(n166), .A2(rt_data[26]), .A3(n192), .A4(rt_data[2]), 
        .Y(n160) );
  AO21X1_LVT U248 ( .A1(n168), .A2(rt_data[10]), .A3(n160), .Y(N479) );
  AO22X1_LVT U249 ( .A1(n166), .A2(rt_data[27]), .A3(n192), .A4(rt_data[3]), 
        .Y(n161) );
  AO21X1_LVT U250 ( .A1(n168), .A2(rt_data[11]), .A3(n161), .Y(N480) );
  AO22X1_LVT U251 ( .A1(n166), .A2(rt_data[28]), .A3(n192), .A4(rt_data[4]), 
        .Y(n162) );
  AO21X1_LVT U252 ( .A1(n168), .A2(rt_data[12]), .A3(n162), .Y(N481) );
  AO22X1_LVT U253 ( .A1(n166), .A2(rt_data[29]), .A3(n192), .A4(rt_data[5]), 
        .Y(n163) );
  AO21X1_LVT U254 ( .A1(n168), .A2(rt_data[13]), .A3(n163), .Y(N482) );
  AO22X1_LVT U255 ( .A1(n166), .A2(rt_data[30]), .A3(n192), .A4(rt_data[6]), 
        .Y(n164) );
  AO21X1_LVT U256 ( .A1(n168), .A2(rt_data[14]), .A3(n164), .Y(N483) );
  AO22X1_LVT U257 ( .A1(n166), .A2(rt_data[31]), .A3(n192), .A4(rt_data[7]), 
        .Y(n167) );
  AO21X1_LVT U258 ( .A1(n168), .A2(rt_data[15]), .A3(n167), .Y(N484) );
  AND2X1_LVT U259 ( .A1(mem_addr_i[0]), .A2(N420), .Y(N421) );
  AND2X1_LVT U263 ( .A1(mem_addr_i[2]), .A2(n170), .Y(N423) );
  AND2X1_LVT U264 ( .A1(mem_addr_i[3]), .A2(n170), .Y(N424) );
  AND2X1_LVT U265 ( .A1(mem_addr_i[4]), .A2(n170), .Y(N425) );
  AND2X1_LVT U266 ( .A1(mem_addr_i[5]), .A2(n170), .Y(N426) );
  AND2X1_LVT U267 ( .A1(mem_addr_i[6]), .A2(n170), .Y(N427) );
  AND2X1_LVT U268 ( .A1(mem_addr_i[7]), .A2(n170), .Y(N428) );
  AND2X1_LVT U269 ( .A1(mem_addr_i[8]), .A2(n170), .Y(N429) );
  AND2X1_LVT U270 ( .A1(mem_addr_i[9]), .A2(n170), .Y(N430) );
  AND2X1_LVT U271 ( .A1(mem_addr_i[10]), .A2(n170), .Y(N431) );
  AND2X1_LVT U272 ( .A1(mem_addr_i[11]), .A2(n170), .Y(N432) );
  AND2X1_LVT U273 ( .A1(mem_addr_i[12]), .A2(n195), .Y(N433) );
  AND2X1_LVT U274 ( .A1(mem_addr_i[13]), .A2(n170), .Y(N434) );
  AND2X1_LVT U275 ( .A1(mem_addr_i[14]), .A2(n195), .Y(N435) );
  AND2X1_LVT U276 ( .A1(mem_addr_i[15]), .A2(n195), .Y(N436) );
  AND2X1_LVT U277 ( .A1(mem_addr_i[16]), .A2(n195), .Y(N437) );
  AND2X1_LVT U279 ( .A1(mem_addr_i[17]), .A2(n195), .Y(N438) );
  AND2X1_LVT U280 ( .A1(mem_addr_i[18]), .A2(n195), .Y(N439) );
  AND2X1_LVT U281 ( .A1(mem_addr_i[19]), .A2(n195), .Y(N440) );
  AND2X1_LVT U282 ( .A1(mem_addr_i[20]), .A2(n195), .Y(N441) );
  AND2X1_LVT U283 ( .A1(mem_addr_i[21]), .A2(n195), .Y(N442) );
  AND2X1_LVT U284 ( .A1(mem_addr_i[22]), .A2(n195), .Y(N443) );
  AND2X1_LVT U285 ( .A1(mem_addr_i[23]), .A2(n195), .Y(N444) );
  AND2X1_LVT U286 ( .A1(mem_addr_i[24]), .A2(n195), .Y(N445) );
  AND2X1_LVT U287 ( .A1(mem_addr_i[25]), .A2(n195), .Y(N446) );
  AND2X1_LVT U288 ( .A1(mem_addr_i[26]), .A2(n195), .Y(N447) );
  AND2X1_LVT U289 ( .A1(mem_addr_i[27]), .A2(n195), .Y(N448) );
  AND2X1_LVT U290 ( .A1(mem_addr_i[28]), .A2(n195), .Y(N449) );
  AND2X1_LVT U291 ( .A1(mem_addr_i[29]), .A2(n195), .Y(N450) );
  AND2X1_LVT U292 ( .A1(mem_addr_i[30]), .A2(n195), .Y(N451) );
  AND2X1_LVT U293 ( .A1(mem_addr_i[31]), .A2(n195), .Y(N452) );
  NAND2X0_LVT U294 ( .A1(n184), .A2(n172), .Y(N528) );
  NAND2X0_LVT U295 ( .A1(n174), .A2(N528), .Y(stallreq) );
  AND2X2_LVT U260 ( .A1(mem_addr_i[1]), .A2(N420), .Y(N422) );
  OR2X4_LVT U261 ( .A1(N420), .A2(N419), .Y(n170) );
  NAND2X4_LVT U19 ( .A1(n145), .A2(n150), .Y(N420) );
  INVX2_LVT U5 ( .A(rst), .Y(n184) );
  INVX1_LVT U9 ( .A(aluop[0]), .Y(n185) );
  INVX1_LVT U10 ( .A(aluop[1]), .Y(n186) );
  INVX1_LVT U20 ( .A(mem_addr_i[0]), .Y(n187) );
  INVX1_LVT U23 ( .A(mem_addr_i[1]), .Y(n188) );
  INVX4_LVT U24 ( .A(n20), .Y(n189) );
  NBUFFX8_LVT U25 ( .A(n4), .Y(n190) );
  NBUFFX8_LVT U26 ( .A(n4), .Y(n191) );
  INVX2_LVT U34 ( .A(n150), .Y(n192) );
  NAND3X2_LVT U33 ( .A1(n184), .A2(n15), .A3(n10), .Y(n11) );
  AO21X2_LVT U56 ( .A1(n119), .A2(n109), .A3(n116), .Y(n131) );
  LATCHX2_LVT \mem_addr_o_reg[0]  ( .CLK(n190), .D(N421), .Q(mem_addr_o[0]) );
  NBUFFX4_LVT U35 ( .A(n131), .Y(n194) );
  NAND3X0_LVT U36 ( .A1(n71), .A2(n119), .A3(n61), .Y(n193) );
  NBUFFX4_LVT U37 ( .A(n170), .Y(n195) );
  NBUFFX4_LVT U38 ( .A(n11), .Y(n196) );
endmodule


module pipe_mem_wb ( clk, rst, mem_reg_waddr, mem_we, mem_reg_wdata, stall, 
        wb_reg_waddr, wb_we, wb_reg_wdata );
  input [4:0] mem_reg_waddr;
  input [31:0] mem_reg_wdata;
  input [5:0] stall;
  output [4:0] wb_reg_waddr;
  output [31:0] wb_reg_wdata;
  input clk, rst, mem_we;
  output wb_we;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n1, n48;

  DFFX1_LVT \wb_reg_wdata_reg[11]  ( .D(n13), .CLK(clk), .Q(wb_reg_wdata[11])
         );
  DFFX1_LVT \wb_reg_wdata_reg[7]  ( .D(n9), .CLK(clk), .Q(wb_reg_wdata[7]) );
  DFFX1_LVT \wb_reg_wdata_reg[6]  ( .D(n8), .CLK(clk), .Q(wb_reg_wdata[6]) );
  DFFX1_LVT wb_we_reg ( .D(n34), .CLK(clk), .Q(wb_we) );
  DFFX1_LVT \wb_reg_waddr_reg[3]  ( .D(n38), .CLK(clk), .Q(wb_reg_waddr[3]) );
  DFFX1_LVT \wb_reg_waddr_reg[4]  ( .D(n39), .CLK(clk), .Q(wb_reg_waddr[4]) );
  DFFX1_LVT \wb_reg_waddr_reg[0]  ( .D(n35), .CLK(clk), .Q(wb_reg_waddr[0]) );
  DFFX1_LVT \wb_reg_waddr_reg[1]  ( .D(n36), .CLK(clk), .Q(wb_reg_waddr[1]) );
  AND2X1_LVT U6 ( .A1(n48), .A2(mem_reg_waddr[4]), .Y(n39) );
  AND2X1_LVT U7 ( .A1(n48), .A2(mem_reg_waddr[3]), .Y(n38) );
  AND2X1_LVT U8 ( .A1(n48), .A2(mem_reg_waddr[2]), .Y(n37) );
  AND2X1_LVT U9 ( .A1(n48), .A2(mem_reg_waddr[1]), .Y(n36) );
  AND2X1_LVT U10 ( .A1(n48), .A2(mem_reg_waddr[0]), .Y(n35) );
  AND2X1_LVT U11 ( .A1(n48), .A2(mem_we), .Y(n34) );
  AND2X1_LVT U12 ( .A1(n48), .A2(mem_reg_wdata[31]), .Y(n33) );
  AND2X1_LVT U13 ( .A1(n48), .A2(mem_reg_wdata[30]), .Y(n32) );
  AND2X1_LVT U14 ( .A1(n48), .A2(mem_reg_wdata[29]), .Y(n31) );
  AND2X1_LVT U15 ( .A1(n48), .A2(mem_reg_wdata[28]), .Y(n30) );
  AND2X1_LVT U16 ( .A1(n48), .A2(mem_reg_wdata[27]), .Y(n29) );
  AND2X1_LVT U17 ( .A1(n48), .A2(mem_reg_wdata[26]), .Y(n28) );
  AND2X1_LVT U18 ( .A1(n48), .A2(mem_reg_wdata[25]), .Y(n27) );
  AND2X1_LVT U19 ( .A1(n48), .A2(mem_reg_wdata[24]), .Y(n26) );
  AND2X1_LVT U20 ( .A1(n48), .A2(mem_reg_wdata[23]), .Y(n25) );
  AND2X1_LVT U22 ( .A1(n48), .A2(mem_reg_wdata[22]), .Y(n24) );
  AND2X1_LVT U23 ( .A1(n1), .A2(mem_reg_wdata[21]), .Y(n23) );
  AND2X1_LVT U24 ( .A1(n48), .A2(mem_reg_wdata[20]), .Y(n22) );
  AND2X1_LVT U25 ( .A1(n48), .A2(mem_reg_wdata[19]), .Y(n21) );
  AND2X1_LVT U26 ( .A1(n48), .A2(mem_reg_wdata[18]), .Y(n20) );
  AND2X1_LVT U27 ( .A1(n48), .A2(mem_reg_wdata[17]), .Y(n19) );
  AND2X1_LVT U28 ( .A1(n48), .A2(mem_reg_wdata[16]), .Y(n18) );
  AND2X1_LVT U29 ( .A1(n48), .A2(mem_reg_wdata[15]), .Y(n17) );
  AND2X1_LVT U30 ( .A1(n48), .A2(mem_reg_wdata[14]), .Y(n16) );
  AND2X1_LVT U31 ( .A1(n48), .A2(mem_reg_wdata[13]), .Y(n15) );
  AND2X1_LVT U32 ( .A1(n48), .A2(mem_reg_wdata[12]), .Y(n14) );
  AND2X1_LVT U33 ( .A1(n48), .A2(mem_reg_wdata[11]), .Y(n13) );
  AND2X1_LVT U34 ( .A1(n48), .A2(mem_reg_wdata[10]), .Y(n12) );
  AND2X1_LVT U35 ( .A1(n48), .A2(mem_reg_wdata[9]), .Y(n11) );
  AND2X1_LVT U36 ( .A1(n48), .A2(mem_reg_wdata[8]), .Y(n10) );
  AND2X1_LVT U38 ( .A1(n48), .A2(mem_reg_wdata[7]), .Y(n9) );
  AND2X1_LVT U39 ( .A1(n48), .A2(mem_reg_wdata[6]), .Y(n8) );
  AND2X1_LVT U40 ( .A1(n48), .A2(mem_reg_wdata[5]), .Y(n7) );
  AND2X1_LVT U41 ( .A1(n48), .A2(mem_reg_wdata[4]), .Y(n6) );
  AND2X1_LVT U42 ( .A1(n48), .A2(mem_reg_wdata[3]), .Y(n5) );
  AND2X1_LVT U43 ( .A1(n48), .A2(mem_reg_wdata[2]), .Y(n4) );
  AND2X1_LVT U44 ( .A1(n48), .A2(mem_reg_wdata[1]), .Y(n3) );
  AND2X1_LVT U45 ( .A1(n48), .A2(mem_reg_wdata[0]), .Y(n2) );
  DFFX2_LVT \wb_reg_wdata_reg[26]  ( .D(n28), .CLK(clk), .Q(wb_reg_wdata[26])
         );
  DFFX2_LVT \wb_reg_wdata_reg[30]  ( .D(n32), .CLK(clk), .Q(wb_reg_wdata[30])
         );
  DFFX2_LVT \wb_reg_wdata_reg[28]  ( .D(n30), .CLK(clk), .Q(wb_reg_wdata[28])
         );
  DFFX2_LVT \wb_reg_wdata_reg[13]  ( .D(n15), .CLK(clk), .Q(wb_reg_wdata[13])
         );
  DFFX2_LVT \wb_reg_wdata_reg[27]  ( .D(n29), .CLK(clk), .Q(wb_reg_wdata[27])
         );
  DFFX2_LVT \wb_reg_wdata_reg[10]  ( .D(n12), .CLK(clk), .Q(wb_reg_wdata[10])
         );
  DFFX2_LVT \wb_reg_wdata_reg[31]  ( .D(n33), .CLK(clk), .Q(wb_reg_wdata[31])
         );
  DFFX2_LVT \wb_reg_wdata_reg[12]  ( .D(n14), .CLK(clk), .Q(wb_reg_wdata[12])
         );
  DFFX2_LVT \wb_reg_wdata_reg[25]  ( .D(n27), .CLK(clk), .Q(wb_reg_wdata[25])
         );
  DFFX2_LVT \wb_reg_wdata_reg[29]  ( .D(n31), .CLK(clk), .Q(wb_reg_wdata[29])
         );
  DFFX2_LVT \wb_reg_wdata_reg[9]  ( .D(n11), .CLK(clk), .Q(wb_reg_wdata[9]) );
  DFFX2_LVT \wb_reg_wdata_reg[14]  ( .D(n16), .CLK(clk), .Q(wb_reg_wdata[14])
         );
  DFFX2_LVT \wb_reg_wdata_reg[16]  ( .D(n18), .CLK(clk), .Q(wb_reg_wdata[16])
         );
  DFFX2_LVT \wb_reg_wdata_reg[15]  ( .D(n17), .CLK(clk), .Q(wb_reg_wdata[15])
         );
  DFFX2_LVT \wb_reg_wdata_reg[23]  ( .D(n25), .CLK(clk), .Q(wb_reg_wdata[23])
         );
  DFFX2_LVT \wb_reg_wdata_reg[19]  ( .D(n21), .CLK(clk), .Q(wb_reg_wdata[19])
         );
  DFFX2_LVT \wb_reg_wdata_reg[20]  ( .D(n22), .CLK(clk), .Q(wb_reg_wdata[20])
         );
  DFFX2_LVT \wb_reg_wdata_reg[24]  ( .D(n26), .CLK(clk), .Q(wb_reg_wdata[24])
         );
  DFFX2_LVT \wb_reg_wdata_reg[18]  ( .D(n20), .CLK(clk), .Q(wb_reg_wdata[18])
         );
  DFFX2_LVT \wb_reg_wdata_reg[22]  ( .D(n24), .CLK(clk), .Q(wb_reg_wdata[22])
         );
  DFFX2_LVT \wb_reg_wdata_reg[8]  ( .D(n10), .CLK(clk), .Q(wb_reg_wdata[8]) );
  DFFX2_LVT \wb_reg_wdata_reg[17]  ( .D(n19), .CLK(clk), .Q(wb_reg_wdata[17])
         );
  DFFX2_LVT \wb_reg_wdata_reg[5]  ( .D(n7), .CLK(clk), .Q(wb_reg_wdata[5]) );
  DFFX2_LVT \wb_reg_wdata_reg[21]  ( .D(n23), .CLK(clk), .Q(wb_reg_wdata[21])
         );
  DFFX2_LVT \wb_reg_wdata_reg[0]  ( .D(n2), .CLK(clk), .Q(wb_reg_wdata[0]) );
  DFFX2_LVT \wb_reg_wdata_reg[1]  ( .D(n3), .CLK(clk), .Q(wb_reg_wdata[1]) );
  DFFX1_LVT \wb_reg_wdata_reg[4]  ( .D(n6), .CLK(clk), .Q(wb_reg_wdata[4]) );
  DFFX1_LVT \wb_reg_wdata_reg[3]  ( .D(n5), .CLK(clk), .Q(wb_reg_wdata[3]) );
  DFFX1_LVT \wb_reg_wdata_reg[2]  ( .D(n4), .CLK(clk), .Q(wb_reg_wdata[2]) );
  DFFX1_LVT \wb_reg_waddr_reg[2]  ( .D(n37), .CLK(clk), .Q(wb_reg_waddr[2]) );
  NOR2X2_LVT U3 ( .A1(stall[4]), .A2(rst), .Y(n1) );
  NBUFFX8_LVT U4 ( .A(n1), .Y(n48) );
endmodule


module riscv_cpu ( clk, rst, mem_data_i, mem_busy_i, mem_done_i, mem_rwe_o, 
        mem_addr_o, mem_sel_o, mem_data_o );
  input [31:0] mem_data_i;
  input [1:0] mem_busy_i;
  input [1:0] mem_done_i;
  output [3:0] mem_rwe_o;
  output [31:0] mem_addr_o;
  output [7:0] mem_sel_o;
  output [31:0] mem_data_o;
  input clk, rst;
  wire   stallreq_if, stallreq_id, stallreq_mem, br, right_one, ex_we_o,
         mem_we_o, id_re1, id_re2, id_we, wb_we, ex_we_i, mem_we_i, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135;
  wire   [5:0] stall;
  wire   [31:0] br_addr;
  wire   [31:0] pc;
  wire   [31:0] if_pc;
  wire   [31:0] if_inst;
  wire   [31:0] id_pc;
  wire   [31:0] id_inst;
  wire   [31:0] id_reg_data1;
  wire   [31:0] id_reg_data2;
  wire   [7:0] ex_aluop;
  wire   [4:0] ex_reg_waddr_o;
  wire   [31:0] ex_reg_wdata;
  wire   [4:0] mem_reg_waddr_o;
  wire   [31:0] mem_reg_wdata_o;
  wire   [4:0] id_reg_addr1;
  wire   [4:0] id_reg_addr2;
  wire   [7:0] id_aluop;
  wire   [2:0] id_alusel;
  wire   [31:0] id_opv1;
  wire   [31:0] id_opv2;
  wire   [4:0] id_reg_waddr;
  wire   [31:0] id_link_addr;
  wire   [31:0] id_mem_offset;
  wire   [4:0] wb_reg_waddr;
  wire   [31:0] wb_reg_wdata;
  wire   [2:0] ex_alusel;
  wire   [31:0] ex_opv1;
  wire   [31:0] ex_opv2;
  wire   [4:0] ex_reg_waddr_i;
  wire   [31:0] ex_link_addr;
  wire   [31:0] ex_mem_offset;
  wire   [31:0] ex_mem_addr;
  wire   [7:0] ex_aluop_o;
  wire   [31:0] ex_rt_data;
  wire   [4:0] mem_reg_waddr_i;
  wire   [31:0] mem_reg_wdata_i;
  wire   [31:0] mem_mem_addr;
  wire   [7:0] mem_aluop;
  wire   [31:0] mem_rt_data;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12;

  stall_ctrl stall_ctrl0 ( .rst(rst), .stallreq_if(stallreq_if), .stallreq_id(
        stallreq_id), .stallreq_ex(1'b0), .stallreq_mem(stallreq_mem), .stall(
        {SYNOPSYS_UNCONNECTED__0, stall[4:0]}) );
  program_counter program_counter0 ( .clk(clk), .rst(rst), .stall({1'b0, 
        stall[4:0]}), .br(br), .br_addr(br_addr), .pc_o(pc), .right_one_o(
        right_one) );
  inst_fetch inst_fetch0 ( .rst(rst), .pc_i(pc), .mem_data_i(mem_data_i), 
        .mem_busy(mem_busy_i), .mem_done(mem_done_i), .br(br), .right_one(
        right_one), .mem_addr_o({n64, n62, n60, n58, n56, n54, n52, n50, n48, 
        n46, n44, n42, n40, n38, n36, n34, n32, n30, n28, n26, n24, n22, n20, 
        n18, n16, n14, n12, n10, n8, n6, n4, n2}), .pc_o(if_pc), .inst_o(
        if_inst), .stallreq(stallreq_if) );
  pipe_if_id pipe_if_id0 ( .clk(clk), .rst(rst), .if_pc(if_pc), .if_inst(
        if_inst), .stall({1'b0, stall[4:0]}), .br(br), .id_pc(id_pc), 
        .id_inst(id_inst) );
  inst_decoder inst_decoder0 ( .rst(rst), .pc({n106, id_pc[30:29], n105, 
        id_pc[27], n104, id_pc[25:24], n103, id_pc[22:4], n102, n101, 
        id_pc[1:0]}), .inst({n100, id_inst[30:4], n99, id_inst[2:0]}), 
        .reg_data1(id_reg_data1), .reg_data2(id_reg_data2), .ex_aluop({1'b0, 
        1'b0, 1'b0, ex_aluop[4:0]}), .ex_we(ex_we_o), .ex_reg_wdata({
        ex_reg_wdata[31:28], n112, n113, ex_reg_wdata[25:20], n116, n117, 
        ex_reg_wdata[17:16], n120, ex_reg_wdata[14:8], n111, ex_reg_wdata[6:3], 
        n118, ex_reg_wdata[1], n119}), .ex_reg_waddr(ex_reg_waddr_o), .mem_we(
        mem_we_o), .mem_reg_wdata(mem_reg_wdata_o), .mem_reg_waddr(
        mem_reg_waddr_o), .re1(id_re1), .re2(id_re2), .reg_addr1(id_reg_addr1), 
        .reg_addr2(id_reg_addr2), .aluop({SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, id_aluop[4:0]}), 
        .alusel(id_alusel), .opv1(id_opv1), .opv2(id_opv2), .reg_waddr(
        id_reg_waddr), .we(id_we), .stallreq(stallreq_id), .br(br), .br_addr(
        br_addr), .link_addr(id_link_addr), .mem_offset(id_mem_offset) );
  regfile regfile0 ( .clk(clk), .rst(rst), .we(wb_we), .waddr(wb_reg_waddr), 
        .wdata({n114, n127, wb_reg_wdata[29:28], n130, wb_reg_wdata[26], n129, 
        wb_reg_wdata[24:22], n132, wb_reg_wdata[20:18], n134, n125, 
        wb_reg_wdata[15:13], n123, n109, wb_reg_wdata[10], n122, n135, n108, 
        n107, n133, n131, n128, n121, n124, n126}), .re1(id_re1), .raddr1(
        id_reg_addr1), .rdata1(id_reg_data1), .re2(id_re2), .raddr2(
        id_reg_addr2), .rdata2(id_reg_data2) );
  pipe_id_ex pipe_id_ex0 ( .clk(clk), .rst(rst), .id_aluop({1'b0, 1'b0, 1'b0, 
        id_aluop[4:0]}), .id_alusel(id_alusel), .id_opv1(id_opv1), .id_opv2(
        id_opv2), .id_reg_waddr(id_reg_waddr), .id_we(id_we), .stall({1'b0, 
        stall[4:0]}), .id_link_addr(id_link_addr), .id_mem_offset(
        id_mem_offset), .ex_aluop({SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, ex_aluop[4:0]}), 
        .ex_alusel(ex_alusel), .ex_opv1(ex_opv1), .ex_opv2(ex_opv2), 
        .ex_reg_waddr(ex_reg_waddr_i), .ex_we(ex_we_i), .ex_link_addr(
        ex_link_addr), .ex_mem_offset(ex_mem_offset) );
  execute_alu execute_alu0 ( .rst(rst), .aluop({1'b0, 1'b0, 1'b0, 
        ex_aluop[4:0]}), .alusel(ex_alusel), .opv1({ex_opv1[31:30], n115, 
        ex_opv1[28:2], n110, n68}), .opv2({n97, n96, n95, n94, n91, n93, n92, 
        n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, n77, 
        n76, ex_opv2[9], n75, n74, n73, n72, n71, n70, n69, n67, n66}), 
        .reg_waddr_i(ex_reg_waddr_i), .we_i(ex_we_i), .link_addr(ex_link_addr), 
        .mem_offset(ex_mem_offset), .reg_waddr_o(ex_reg_waddr_o), .we_o(
        ex_we_o), .reg_wdata(ex_reg_wdata), .mem_addr(ex_mem_addr), .ex_aluop(
        {SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, ex_aluop_o[4:0]}), .rt_data(ex_rt_data) );
  pipe_ex_mem pipe_ex_mem0 ( .clk(clk), .rst(rst), .ex_reg_waddr(
        ex_reg_waddr_o), .ex_we(ex_we_o), .ex_reg_wdata({ex_reg_wdata[31:28], 
        n112, n113, ex_reg_wdata[25:20], n116, n117, ex_reg_wdata[17:16], n120, 
        ex_reg_wdata[14:3], n118, ex_reg_wdata[1], n119}), .stall({1'b0, 
        stall[4:0]}), .ex_mem_addr(ex_mem_addr), .ex_aluop({1'b0, 1'b0, 1'b0, 
        ex_aluop_o[4:0]}), .ex_rt_data(ex_rt_data), .mem_reg_waddr(
        mem_reg_waddr_i), .mem_we(mem_we_i), .mem_reg_wdata(mem_reg_wdata_i), 
        .mem_mem_addr(mem_mem_addr), .mem_aluop({SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, mem_aluop[4:0]}), 
        .mem_rt_data(mem_rt_data) );
  stage_mem stage_mem0 ( .rst(rst), .reg_waddr_i(mem_reg_waddr_i), .we_i(
        mem_we_i), .reg_wdata_i(mem_reg_wdata_i), .mem_addr_i({
        mem_mem_addr[31:1], n98}), .aluop({1'b0, 1'b0, 1'b0, mem_aluop[4:0]}), 
        .rt_data(mem_rt_data), .mem_data_i(mem_data_i), .mem_busy(mem_busy_i), 
        .mem_done(mem_done_i), .reg_waddr_o(mem_reg_waddr_o), .we_o(mem_we_o), 
        .reg_wdata_o(mem_reg_wdata_o), .mem_addr_o({n65, n63, n61, n59, n57, 
        n55, n53, n51, n49, n47, n45, n43, n41, n39, n37, n35, n33, n31, n29, 
        n27, n25, n23, n21, n19, n17, n15, n13, n11, n9, n7, n5, n3}), 
        .mem_data_o(mem_data_o), .stallreq(stallreq_mem) );
  pipe_mem_wb pipe_mem_wb0 ( .clk(clk), .rst(rst), .mem_reg_waddr(
        mem_reg_waddr_o), .mem_we(mem_we_o), .mem_reg_wdata(mem_reg_wdata_o), 
        .stall({1'b0, stall[4:0]}), .wb_reg_waddr(wb_reg_waddr), .wb_we(wb_we), 
        .wb_reg_wdata(wb_reg_wdata) );
  AND2X1_LVT U3 ( .A1(n2), .A2(n3), .Y(mem_addr_o[0]) );
  AND2X1_LVT U4 ( .A1(n4), .A2(n5), .Y(mem_addr_o[1]) );
  AND2X1_LVT U5 ( .A1(n6), .A2(n7), .Y(mem_addr_o[2]) );
  AND2X1_LVT U6 ( .A1(n8), .A2(n9), .Y(mem_addr_o[3]) );
  AND2X1_LVT U7 ( .A1(n10), .A2(n11), .Y(mem_addr_o[4]) );
  AND2X1_LVT U8 ( .A1(n12), .A2(n13), .Y(mem_addr_o[5]) );
  AND2X1_LVT U9 ( .A1(n14), .A2(n15), .Y(mem_addr_o[6]) );
  AND2X1_LVT U10 ( .A1(n16), .A2(n17), .Y(mem_addr_o[7]) );
  AND2X1_LVT U11 ( .A1(n18), .A2(n19), .Y(mem_addr_o[8]) );
  AND2X1_LVT U12 ( .A1(n20), .A2(n21), .Y(mem_addr_o[9]) );
  AND2X1_LVT U13 ( .A1(n22), .A2(n23), .Y(mem_addr_o[10]) );
  AND2X1_LVT U14 ( .A1(n24), .A2(n25), .Y(mem_addr_o[11]) );
  AND2X1_LVT U15 ( .A1(n26), .A2(n27), .Y(mem_addr_o[12]) );
  AND2X1_LVT U16 ( .A1(n28), .A2(n29), .Y(mem_addr_o[13]) );
  AND2X1_LVT U17 ( .A1(n30), .A2(n31), .Y(mem_addr_o[14]) );
  AND2X1_LVT U18 ( .A1(n32), .A2(n33), .Y(mem_addr_o[15]) );
  AND2X1_LVT U19 ( .A1(n34), .A2(n35), .Y(mem_addr_o[16]) );
  AND2X1_LVT U20 ( .A1(n36), .A2(n37), .Y(mem_addr_o[17]) );
  AND2X1_LVT U21 ( .A1(n38), .A2(n39), .Y(mem_addr_o[18]) );
  AND2X1_LVT U22 ( .A1(n40), .A2(n41), .Y(mem_addr_o[19]) );
  AND2X1_LVT U23 ( .A1(n42), .A2(n43), .Y(mem_addr_o[20]) );
  AND2X1_LVT U24 ( .A1(n44), .A2(n45), .Y(mem_addr_o[21]) );
  AND2X1_LVT U25 ( .A1(n46), .A2(n47), .Y(mem_addr_o[22]) );
  AND2X1_LVT U26 ( .A1(n48), .A2(n49), .Y(mem_addr_o[23]) );
  AND2X1_LVT U27 ( .A1(n50), .A2(n51), .Y(mem_addr_o[24]) );
  AND2X1_LVT U28 ( .A1(n52), .A2(n53), .Y(mem_addr_o[25]) );
  AND2X1_LVT U29 ( .A1(n54), .A2(n55), .Y(mem_addr_o[26]) );
  AND2X1_LVT U30 ( .A1(n56), .A2(n57), .Y(mem_addr_o[27]) );
  AND2X1_LVT U31 ( .A1(n58), .A2(n59), .Y(mem_addr_o[28]) );
  AND2X1_LVT U32 ( .A1(n60), .A2(n61), .Y(mem_addr_o[29]) );
  AND2X1_LVT U33 ( .A1(n62), .A2(n63), .Y(mem_addr_o[30]) );
  AND2X1_LVT U34 ( .A1(n64), .A2(n65), .Y(mem_addr_o[31]) );
  NBUFFX4_LVT U35 ( .A(ex_opv2[0]), .Y(n66) );
  NBUFFX4_LVT U36 ( .A(ex_opv2[1]), .Y(n67) );
  NBUFFX4_LVT U37 ( .A(ex_opv1[0]), .Y(n68) );
  NBUFFX4_LVT U38 ( .A(ex_opv2[2]), .Y(n69) );
  NBUFFX4_LVT U39 ( .A(ex_opv2[3]), .Y(n70) );
  NBUFFX4_LVT U40 ( .A(ex_opv2[4]), .Y(n71) );
  NBUFFX4_LVT U41 ( .A(ex_opv2[5]), .Y(n72) );
  NBUFFX4_LVT U42 ( .A(ex_opv2[6]), .Y(n73) );
  NBUFFX4_LVT U43 ( .A(ex_opv2[7]), .Y(n74) );
  NBUFFX4_LVT U44 ( .A(ex_opv2[8]), .Y(n75) );
  NBUFFX4_LVT U45 ( .A(ex_opv2[10]), .Y(n76) );
  NBUFFX4_LVT U46 ( .A(ex_opv2[11]), .Y(n77) );
  NBUFFX4_LVT U47 ( .A(ex_opv2[12]), .Y(n78) );
  NBUFFX4_LVT U48 ( .A(ex_opv2[13]), .Y(n79) );
  NBUFFX4_LVT U49 ( .A(ex_opv2[14]), .Y(n80) );
  NBUFFX4_LVT U50 ( .A(ex_opv2[15]), .Y(n81) );
  NBUFFX4_LVT U51 ( .A(ex_opv2[16]), .Y(n82) );
  NBUFFX4_LVT U52 ( .A(ex_opv2[17]), .Y(n83) );
  NBUFFX4_LVT U53 ( .A(ex_opv2[18]), .Y(n84) );
  NBUFFX4_LVT U54 ( .A(ex_opv2[19]), .Y(n85) );
  NBUFFX4_LVT U55 ( .A(ex_opv2[20]), .Y(n86) );
  NBUFFX4_LVT U56 ( .A(ex_opv2[21]), .Y(n87) );
  NBUFFX4_LVT U57 ( .A(ex_opv2[22]), .Y(n88) );
  NBUFFX4_LVT U58 ( .A(ex_opv2[23]), .Y(n89) );
  NBUFFX4_LVT U59 ( .A(ex_opv2[24]), .Y(n90) );
  NBUFFX4_LVT U60 ( .A(ex_opv2[27]), .Y(n91) );
  NBUFFX4_LVT U61 ( .A(ex_opv2[25]), .Y(n92) );
  NBUFFX4_LVT U62 ( .A(ex_opv2[26]), .Y(n93) );
  NBUFFX4_LVT U63 ( .A(ex_opv2[28]), .Y(n94) );
  NBUFFX4_LVT U64 ( .A(ex_opv2[29]), .Y(n95) );
  NBUFFX4_LVT U65 ( .A(ex_opv2[30]), .Y(n96) );
  NBUFFX4_LVT U66 ( .A(ex_opv2[31]), .Y(n97) );
  NBUFFX4_LVT U67 ( .A(mem_mem_addr[0]), .Y(n98) );
  NBUFFX4_LVT U68 ( .A(id_inst[3]), .Y(n99) );
  NBUFFX4_LVT U69 ( .A(id_inst[31]), .Y(n100) );
  NBUFFX4_LVT U70 ( .A(id_pc[2]), .Y(n101) );
  NBUFFX4_LVT U71 ( .A(id_pc[3]), .Y(n102) );
  NBUFFX4_LVT U72 ( .A(id_pc[23]), .Y(n103) );
  NBUFFX4_LVT U73 ( .A(id_pc[26]), .Y(n104) );
  NBUFFX4_LVT U74 ( .A(id_pc[28]), .Y(n105) );
  NBUFFX4_LVT U75 ( .A(id_pc[31]), .Y(n106) );
  NBUFFX8_LVT U76 ( .A(wb_reg_wdata[6]), .Y(n107) );
  NBUFFX8_LVT U77 ( .A(wb_reg_wdata[7]), .Y(n108) );
  NBUFFX8_LVT U78 ( .A(wb_reg_wdata[11]), .Y(n109) );
  NBUFFX4_LVT U79 ( .A(ex_opv1[1]), .Y(n110) );
  NBUFFX4_LVT U80 ( .A(ex_reg_wdata[7]), .Y(n111) );
  NBUFFX4_LVT U81 ( .A(ex_reg_wdata[27]), .Y(n112) );
  NBUFFX4_LVT U82 ( .A(ex_reg_wdata[26]), .Y(n113) );
  NBUFFX4_LVT U83 ( .A(wb_reg_wdata[31]), .Y(n114) );
  NBUFFX4_LVT U84 ( .A(ex_opv1[29]), .Y(n115) );
  NBUFFX8_LVT U85 ( .A(wb_reg_wdata[16]), .Y(n125) );
  NBUFFX8_LVT U86 ( .A(wb_reg_wdata[27]), .Y(n130) );
  NBUFFX8_LVT U87 ( .A(wb_reg_wdata[25]), .Y(n129) );
  NBUFFX8_LVT U88 ( .A(wb_reg_wdata[9]), .Y(n122) );
  NBUFFX8_LVT U89 ( .A(wb_reg_wdata[12]), .Y(n123) );
  NBUFFX8_LVT U90 ( .A(wb_reg_wdata[30]), .Y(n127) );
  NBUFFX4_LVT U91 ( .A(ex_reg_wdata[19]), .Y(n116) );
  NBUFFX4_LVT U92 ( .A(ex_reg_wdata[18]), .Y(n117) );
  NBUFFX4_LVT U93 ( .A(ex_reg_wdata[2]), .Y(n118) );
  NBUFFX4_LVT U94 ( .A(ex_reg_wdata[0]), .Y(n119) );
  NBUFFX4_LVT U95 ( .A(ex_reg_wdata[15]), .Y(n120) );
  NBUFFX8_LVT U96 ( .A(wb_reg_wdata[2]), .Y(n121) );
  NBUFFX8_LVT U97 ( .A(wb_reg_wdata[1]), .Y(n124) );
  NBUFFX8_LVT U98 ( .A(wb_reg_wdata[0]), .Y(n126) );
  NBUFFX8_LVT U99 ( .A(wb_reg_wdata[3]), .Y(n128) );
  NBUFFX8_LVT U100 ( .A(wb_reg_wdata[4]), .Y(n131) );
  NBUFFX8_LVT U101 ( .A(wb_reg_wdata[21]), .Y(n132) );
  NBUFFX8_LVT U102 ( .A(wb_reg_wdata[5]), .Y(n133) );
  NBUFFX8_LVT U103 ( .A(wb_reg_wdata[17]), .Y(n134) );
  NBUFFX8_LVT U104 ( .A(wb_reg_wdata[8]), .Y(n135) );
